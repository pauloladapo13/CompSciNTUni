<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-7.65098,9.16148,136.161,-73.3452</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>54.5,-4.5</position>
<gparam>LABEL_TEXT Front Panel</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AI_XOR4</type>
<position>19,-18.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>128 </input>
<input>
<ID>IN_2</ID>251 </input>
<input>
<ID>IN_3</ID>250 </input>
<output>
<ID>OUT</ID>740 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>8.5,-15.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>5,-25</position>
<output>
<ID>OUT_0</ID>250 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>DE_TO</type>
<position>39,-18.5</position>
<input>
<ID>IN_0</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>264</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>71,-33</position>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>273 </input>
<input>
<ID>IN_2</ID>274 </input>
<input>
<ID>IN_3</ID>275 </input>
<input>
<ID>IN_4</ID>276 </input>
<input>
<ID>IN_5</ID>277 </input>
<input>
<ID>IN_6</ID>278 </input>
<input>
<ID>IN_7</ID>279 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>266</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>117.5,-31</position>
<input>
<ID>IN_0</ID>263 </input>
<input>
<ID>IN_1</ID>264 </input>
<input>
<ID>IN_2</ID>266 </input>
<input>
<ID>IN_3</ID>267 </input>
<input>
<ID>IN_4</ID>268 </input>
<input>
<ID>IN_5</ID>269 </input>
<input>
<ID>IN_6</ID>270 </input>
<input>
<ID>IN_7</ID>271 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 35</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>268</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>108,-59.5</position>
<input>
<ID>IN_0</ID>312 </input>
<input>
<ID>IN_1</ID>286 </input>
<input>
<ID>IN_2</ID>285 </input>
<input>
<ID>IN_3</ID>284 </input>
<input>
<ID>IN_4</ID>283 </input>
<input>
<ID>IN_5</ID>282 </input>
<input>
<ID>IN_6</ID>281 </input>
<input>
<ID>IN_7</ID>280 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>270</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>81.5,-61.5</position>
<input>
<ID>IN_0</ID>330 </input>
<input>
<ID>IN_1</ID>316 </input>
<input>
<ID>IN_2</ID>314 </input>
<input>
<ID>IN_3</ID>313 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>272</ID>
<type>AA_TOGGLE</type>
<position>5,-41</position>
<output>
<ID>OUT_0</ID>248 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>274</ID>
<type>DE_TO</type>
<position>14.5,-41</position>
<input>
<ID>IN_0</ID>248 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>662</ID>
<type>GA_LED</type>
<position>107.5,-8</position>
<input>
<ID>N_in0</ID>720 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>278</ID>
<type>DA_FROM</type>
<position>2.5,-21.5</position>
<input>
<ID>IN_0</ID>251 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck3</lparam></gate>
<gate>
<ID>670</ID>
<type>DA_FROM</type>
<position>104,-8</position>
<input>
<ID>IN_0</ID>720 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>672</ID>
<type>GA_LED</type>
<position>107.5,-12</position>
<input>
<ID>N_in0</ID>721 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>674</ID>
<type>DA_FROM</type>
<position>104,-12</position>
<input>
<ID>IN_0</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Execute</lparam></gate>
<gate>
<ID>294</ID>
<type>DA_FROM</type>
<position>53.5,-22.5</position>
<input>
<ID>IN_0</ID>279 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>295</ID>
<type>DA_FROM</type>
<position>54,-25</position>
<input>
<ID>IN_0</ID>278 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>296</ID>
<type>DA_FROM</type>
<position>53.5,-28.5</position>
<input>
<ID>IN_0</ID>277 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>297</ID>
<type>DA_FROM</type>
<position>54,-31</position>
<input>
<ID>IN_0</ID>276 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>298</ID>
<type>DA_FROM</type>
<position>54,-34</position>
<input>
<ID>IN_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>299</ID>
<type>DA_FROM</type>
<position>55,-36.5</position>
<input>
<ID>IN_0</ID>274 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>300</ID>
<type>DA_FROM</type>
<position>54,-40</position>
<input>
<ID>IN_0</ID>273 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>301</ID>
<type>DA_FROM</type>
<position>54.5,-42.5</position>
<input>
<ID>IN_0</ID>272 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>302</ID>
<type>DA_FROM</type>
<position>99.5,-17.5</position>
<input>
<ID>IN_0</ID>271 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>303</ID>
<type>DA_FROM</type>
<position>100,-20</position>
<input>
<ID>IN_0</ID>270 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>304</ID>
<type>DA_FROM</type>
<position>99,-23</position>
<input>
<ID>IN_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>305</ID>
<type>DA_FROM</type>
<position>100,-26</position>
<input>
<ID>IN_0</ID>268 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>306</ID>
<type>DA_FROM</type>
<position>100,-28</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>307</ID>
<type>DA_FROM</type>
<position>100,-31</position>
<input>
<ID>IN_0</ID>266 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>308</ID>
<type>DA_FROM</type>
<position>99.5,-34</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>309</ID>
<type>DA_FROM</type>
<position>99.5,-38</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>312</ID>
<type>DA_FROM</type>
<position>70,-58.5</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 11</lparam></gate>
<gate>
<ID>313</ID>
<type>DA_FROM</type>
<position>70,-61</position>
<input>
<ID>IN_0</ID>314 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 10</lparam></gate>
<gate>
<ID>314</ID>
<type>DA_FROM</type>
<position>70,-63</position>
<input>
<ID>IN_0</ID>316 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 9</lparam></gate>
<gate>
<ID>315</ID>
<type>DA_FROM</type>
<position>70,-65.5</position>
<input>
<ID>IN_0</ID>330 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 8</lparam></gate>
<gate>
<ID>316</ID>
<type>DA_FROM</type>
<position>97,-52</position>
<input>
<ID>IN_0</ID>280 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 7</lparam></gate>
<gate>
<ID>317</ID>
<type>DA_FROM</type>
<position>97,-54.5</position>
<input>
<ID>IN_0</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 6</lparam></gate>
<gate>
<ID>318</ID>
<type>DA_FROM</type>
<position>97,-56.5</position>
<input>
<ID>IN_0</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 5</lparam></gate>
<gate>
<ID>319</ID>
<type>DA_FROM</type>
<position>97,-59</position>
<input>
<ID>IN_0</ID>283 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 4</lparam></gate>
<gate>
<ID>320</ID>
<type>DA_FROM</type>
<position>97,-62</position>
<input>
<ID>IN_0</ID>284 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 3</lparam></gate>
<gate>
<ID>321</ID>
<type>DA_FROM</type>
<position>97,-65</position>
<input>
<ID>IN_0</ID>285 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 2</lparam></gate>
<gate>
<ID>322</ID>
<type>DA_FROM</type>
<position>97,-67</position>
<input>
<ID>IN_0</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 1</lparam></gate>
<gate>
<ID>323</ID>
<type>DA_FROM</type>
<position>97,-69.5</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 0</lparam></gate>
<gate>
<ID>148</ID>
<type>DA_FROM</type>
<position>8,-18.5</position>
<input>
<ID>IN_0</ID>128 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck2</lparam></gate>
<gate>
<ID>746</ID>
<type>BB_CLOCK</type>
<position>5,-29.5</position>
<output>
<ID>CLK</ID>742 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 50</lparam></gate>
<gate>
<ID>753</ID>
<type>AI_XOR2</type>
<position>30.5,-22.5</position>
<input>
<ID>IN_0</ID>740 </input>
<input>
<ID>IN_1</ID>741 </input>
<output>
<ID>OUT</ID>739 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>755</ID>
<type>AA_AND2</type>
<position>19,-30.5</position>
<input>
<ID>IN_0</ID>742 </input>
<input>
<ID>IN_1</ID>743 </input>
<output>
<ID>OUT</ID>741 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>757</ID>
<type>AA_TOGGLE</type>
<position>6.5,-36.5</position>
<output>
<ID>OUT_0</ID>743 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>759</ID>
<type>AA_LABEL</type>
<position>1,-36</position>
<gparam>LABEL_TEXT Run</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10.5,-15.5,16,-15.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-41,12.5,-41</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<connection>
<GID>272</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-25,11.5,-21.5</points>
<intersection>-25 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-21.5,16,-21.5</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-25,11.5,-25</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-21.5,10,-19.5</points>
<intersection>-21.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-19.5,16,-19.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-21.5,10,-21.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,-38,109,-34</points>
<intersection>-38 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109,-34,112.5,-34</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101.5,-38,109,-38</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>109 0</intersection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-34,107,-33</points>
<intersection>-34 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-33,112.5,-33</points>
<connection>
<GID>266</GID>
<name>IN_1</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101.5,-34,107,-34</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-32,107,-31</points>
<intersection>-32 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-32,112.5,-32</points>
<connection>
<GID>266</GID>
<name>IN_2</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102,-31,107,-31</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-31,107.5,-28</points>
<intersection>-31 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-31,112.5,-31</points>
<connection>
<GID>266</GID>
<name>IN_3</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102,-28,107.5,-28</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-30,108.5,-26</points>
<intersection>-30 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-30,112.5,-30</points>
<connection>
<GID>266</GID>
<name>IN_4</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102,-26,108.5,-26</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-29,109.5,-23</points>
<intersection>-29 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-29,112.5,-29</points>
<connection>
<GID>266</GID>
<name>IN_5</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101,-23,109.5,-23</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-28,110,-20</points>
<intersection>-28 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-28,112.5,-28</points>
<connection>
<GID>266</GID>
<name>IN_6</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102,-20,110,-20</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-27,111.5,-17.5</points>
<intersection>-27 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-27,112.5,-27</points>
<connection>
<GID>266</GID>
<name>IN_7</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101.5,-17.5,111.5,-17.5</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-42.5,63,-36</points>
<intersection>-42.5 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-36,66,-36</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-42.5,63,-42.5</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-40,61,-35</points>
<intersection>-40 2</intersection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-35,66,-35</points>
<connection>
<GID>264</GID>
<name>IN_1</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-40,61,-40</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-36.5,60,-34</points>
<intersection>-36.5 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,-34,66,-34</points>
<connection>
<GID>264</GID>
<name>IN_2</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-36.5,60,-36.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-34,61,-33</points>
<intersection>-34 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-33,66,-33</points>
<connection>
<GID>264</GID>
<name>IN_3</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-34,61,-34</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-32,58,-31</points>
<intersection>-32 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-32,66,-32</points>
<connection>
<GID>264</GID>
<name>IN_4</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-31,58,-31</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-31,60.5,-28.5</points>
<intersection>-31 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-31,66,-31</points>
<connection>
<GID>264</GID>
<name>IN_5</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-28.5,60.5,-28.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-30,61,-25</points>
<intersection>-30 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-30,66,-30</points>
<connection>
<GID>264</GID>
<name>IN_6</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-25,61,-25</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-29,62,-22.5</points>
<intersection>-29 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-29,66,-29</points>
<connection>
<GID>264</GID>
<name>IN_7</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-22.5,62,-22.5</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-55.5,102,-52</points>
<intersection>-55.5 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-55.5,103,-55.5</points>
<connection>
<GID>268</GID>
<name>IN_7</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-52,102,-52</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-56.5,101,-54.5</points>
<intersection>-56.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-56.5,103,-56.5</points>
<connection>
<GID>268</GID>
<name>IN_6</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-54.5,101,-54.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-57.5,100,-56.5</points>
<intersection>-57.5 1</intersection>
<intersection>-56.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-57.5,103,-57.5</points>
<connection>
<GID>268</GID>
<name>IN_5</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-56.5,100,-56.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-59,101,-58.5</points>
<intersection>-59 2</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-58.5,103,-58.5</points>
<connection>
<GID>268</GID>
<name>IN_4</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-59,101,-59</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-62,100,-59.5</points>
<intersection>-62 2</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-59.5,103,-59.5</points>
<connection>
<GID>268</GID>
<name>IN_3</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-62,100,-62</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-65,100.5,-60.5</points>
<intersection>-65 2</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-60.5,103,-60.5</points>
<connection>
<GID>268</GID>
<name>IN_2</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-65,100.5,-65</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-67,101,-61.5</points>
<intersection>-67 2</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-61.5,103,-61.5</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-67,101,-67</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-69.5,102,-62.5</points>
<intersection>-69.5 2</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-62.5,103,-62.5</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-69.5,102,-69.5</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-59.5,75,-58.5</points>
<intersection>-59.5 1</intersection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-59.5,78.5,-59.5</points>
<connection>
<GID>270</GID>
<name>IN_3</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-58.5,75,-58.5</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-61,75,-60.5</points>
<intersection>-61 2</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-60.5,78.5,-60.5</points>
<connection>
<GID>270</GID>
<name>IN_2</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-61,75,-61</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-63,75,-61.5</points>
<intersection>-63 2</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-61.5,78.5,-61.5</points>
<connection>
<GID>270</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-63,75,-63</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-17.5,16,-17.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>10 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>10,-18.5,10,-17.5</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>-17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-65.5,75.5,-62.5</points>
<intersection>-65.5 2</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-62.5,78.5,-62.5</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-65.5,75.5,-65.5</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>720</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106,-8,106.5,-8</points>
<connection>
<GID>662</GID>
<name>N_in0</name></connection>
<connection>
<GID>670</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>721</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106,-12,106.5,-12</points>
<connection>
<GID>672</GID>
<name>N_in0</name></connection>
<connection>
<GID>674</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-22.5,35,-18.5</points>
<intersection>-22.5 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-18.5,37,-18.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-22.5,35,-22.5</points>
<connection>
<GID>753</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-21.5,25,-18.5</points>
<intersection>-21.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-21.5,27.5,-21.5</points>
<connection>
<GID>753</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-18.5,25,-18.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>741</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-30.5,24.5,-23.5</points>
<intersection>-30.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-23.5,27.5,-23.5</points>
<connection>
<GID>753</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-30.5,24.5,-30.5</points>
<connection>
<GID>755</GID>
<name>OUT</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>742</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9,-29.5,16,-29.5</points>
<connection>
<GID>755</GID>
<name>IN_0</name></connection>
<connection>
<GID>746</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>743</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-36.5,12,-31.5</points>
<intersection>-36.5 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-31.5,16,-31.5</points>
<connection>
<GID>755</GID>
<name>IN_1</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-36.5,12,-36.5</points>
<connection>
<GID>757</GID>
<name>OUT_0</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>2.50963,5.1965,124.09,-64.5556</PageViewport>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>47.5,-3.5</position>
<gparam>LABEL_TEXT Memory</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AI_RAM_12x16</type>
<position>55,-27</position>
<input>
<ID>ADDRESS_0</ID>19 </input>
<input>
<ID>ADDRESS_1</ID>18 </input>
<input>
<ID>ADDRESS_10</ID>9 </input>
<input>
<ID>ADDRESS_11</ID>8 </input>
<input>
<ID>ADDRESS_2</ID>17 </input>
<input>
<ID>ADDRESS_3</ID>16 </input>
<input>
<ID>ADDRESS_4</ID>15 </input>
<input>
<ID>ADDRESS_5</ID>14 </input>
<input>
<ID>ADDRESS_6</ID>13 </input>
<input>
<ID>ADDRESS_7</ID>12 </input>
<input>
<ID>ADDRESS_8</ID>11 </input>
<input>
<ID>ADDRESS_9</ID>10 </input>
<input>
<ID>DATA_IN_0</ID>28 </input>
<input>
<ID>DATA_IN_1</ID>29 </input>
<input>
<ID>DATA_IN_10</ID>25 </input>
<input>
<ID>DATA_IN_11</ID>24 </input>
<input>
<ID>DATA_IN_12</ID>23 </input>
<input>
<ID>DATA_IN_13</ID>22 </input>
<input>
<ID>DATA_IN_14</ID>21 </input>
<input>
<ID>DATA_IN_15</ID>20 </input>
<input>
<ID>DATA_IN_2</ID>30 </input>
<input>
<ID>DATA_IN_3</ID>31 </input>
<input>
<ID>DATA_IN_4</ID>32 </input>
<input>
<ID>DATA_IN_5</ID>33 </input>
<input>
<ID>DATA_IN_6</ID>34 </input>
<input>
<ID>DATA_IN_7</ID>35 </input>
<input>
<ID>DATA_IN_8</ID>27 </input>
<input>
<ID>DATA_IN_9</ID>26 </input>
<output>
<ID>DATA_OUT_0</ID>28 </output>
<output>
<ID>DATA_OUT_1</ID>29 </output>
<output>
<ID>DATA_OUT_10</ID>25 </output>
<output>
<ID>DATA_OUT_11</ID>24 </output>
<output>
<ID>DATA_OUT_12</ID>23 </output>
<output>
<ID>DATA_OUT_13</ID>22 </output>
<output>
<ID>DATA_OUT_14</ID>21 </output>
<output>
<ID>DATA_OUT_15</ID>20 </output>
<output>
<ID>DATA_OUT_2</ID>30 </output>
<output>
<ID>DATA_OUT_3</ID>31 </output>
<output>
<ID>DATA_OUT_4</ID>32 </output>
<output>
<ID>DATA_OUT_5</ID>33 </output>
<output>
<ID>DATA_OUT_6</ID>34 </output>
<output>
<ID>DATA_OUT_7</ID>35 </output>
<output>
<ID>DATA_OUT_8</ID>27 </output>
<output>
<ID>DATA_OUT_9</ID>26 </output>
<input>
<ID>ENABLE_0</ID>7 </input>
<input>
<ID>write_clock</ID>1 </input>
<input>
<ID>write_enable</ID>6 </input>
<gparam>angle 0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:337 57343</lparam></gate>
<gate>
<ID>8</ID>
<type>DA_FROM</type>
<position>82.5,-25.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>76.5,-28</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Mem Write</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>76.5,-31.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Mem Read</lparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>32.5,-10</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 11</lparam></gate>
<gate>
<ID>27</ID>
<type>DA_FROM</type>
<position>32.5,-12.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 10</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>32.5,-14.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 9</lparam></gate>
<gate>
<ID>29</ID>
<type>DA_FROM</type>
<position>32.5,-17</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 8</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>32.5,-20</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 7</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>32.5,-22.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 6</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>32.5,-24.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 5</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>32.5,-27</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 4</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>32.5,-30</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 3</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>32.5,-33</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 2</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>32.5,-35</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 1</lparam></gate>
<gate>
<ID>37</ID>
<type>DA_FROM</type>
<position>32.5,-37.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 0</lparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>32.5,-41.5</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>32.5,-44.5</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>41</ID>
<type>DE_TO</type>
<position>32,-47.5</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>32,-50.5</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>43</ID>
<type>DE_TO</type>
<position>32,-54</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>32,-57</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>31.5,-60</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>31.5,-63</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>66,-41.5</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>49</ID>
<type>DE_TO</type>
<position>66,-44.5</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>50</ID>
<type>DE_TO</type>
<position>66,-47</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>51</ID>
<type>DE_TO</type>
<position>66,-50</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>52</ID>
<type>DE_TO</type>
<position>66,-53.5</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>53</ID>
<type>DE_TO</type>
<position>66,-56.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>54</ID>
<type>DE_TO</type>
<position>66,-59</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>55</ID>
<type>DE_TO</type>
<position>66,-62</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,-25.5,80.5,-25.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>write_clock</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-28,69,-26.5</points>
<intersection>-28 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-26.5,69,-26.5</points>
<connection>
<GID>6</GID>
<name>write_enable</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-28,74.5,-28</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-31.5,68,-27.5</points>
<intersection>-31.5 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-27.5,68,-27.5</points>
<connection>
<GID>6</GID>
<name>ENABLE_0</name></connection>
<intersection>68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-31.5,74.5,-31.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-10,46,-10</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>46 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>46,-21.5,46,-10</points>
<connection>
<GID>6</GID>
<name>ADDRESS_11</name></connection>
<intersection>-10 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-22.5,45,-12.5</points>
<intersection>-22.5 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-22.5,46,-22.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_10</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-12.5,45,-12.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-23.5,44,-14.5</points>
<intersection>-23.5 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-23.5,46,-23.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_9</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-14.5,44,-14.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-17,43.5,-17</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>43.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43.5,-24.5,43.5,-17</points>
<intersection>-24.5 4</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43.5,-24.5,46,-24.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_8</name></connection>
<intersection>43.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-25.5,40,-20</points>
<intersection>-25.5 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-25.5,46,-25.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_7</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-20,40,-20</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-26.5,46,-26.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_6</name></connection>
<intersection>38 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38,-26.5,38,-22.5</points>
<intersection>-26.5 1</intersection>
<intersection>-22.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>34.5,-22.5,38,-22.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>38 3</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-27.5,37,-24.5</points>
<intersection>-27.5 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-27.5,46,-27.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_5</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-24.5,37,-24.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-28.5,35.5,-27</points>
<intersection>-28.5 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-28.5,46,-28.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_4</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-27,35.5,-27</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-30,40,-29.5</points>
<intersection>-30 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-29.5,46,-29.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_3</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-30,40,-30</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-33,41.5,-30.5</points>
<intersection>-33 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-30.5,46,-30.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_2</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-33,41.5,-33</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-35,43,-31.5</points>
<intersection>-35 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-31.5,46,-31.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_1</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-35,43,-35</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-37.5,45,-32.5</points>
<intersection>-37.5 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-32.5,46,-32.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-37.5,45,-37.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-41.5,47.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_15</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_15</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-41.5,47.5,-41.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-44.5,48.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_14</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_14</name></connection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-44.5,48.5,-44.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-47.5,49.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_13</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_13</name></connection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-47.5,49.5,-47.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-50.5,50.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_12</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_12</name></connection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-50.5,50.5,-50.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-54,51.5,-54</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>51.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>51.5,-54,51.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_11</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_11</name></connection>
<intersection>-54 1</intersection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-57,52.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_10</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_10</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-57,52.5,-57</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-60,53.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_9</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_9</name></connection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-60,53.5,-60</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-63,54.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_8</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_8</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-63,54.5,-63</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-41.5,62.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_0</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-41.5,64,-41.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-44.5,61.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_1</name></connection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-44.5,64,-44.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-47,60.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_2</name></connection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-47,64,-47</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-50,59.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_3</name></connection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-50,64,-50</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-53.5,58.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_4</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-53.5,64,-53.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-56.5,57.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_5</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-56.5,64,-56.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-59,56.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_6</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-59,64,-59</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-62,55.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_7</name></connection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-62,64,-62</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-88.0328,65.7758,200.158,-99.5627</PageViewport>
<gate>
<ID>772</ID>
<type>DE_TO</type>
<position>104.5,-68</position>
<input>
<ID>IN_0</ID>681 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I1</lparam></gate>
<gate>
<ID>773</ID>
<type>DE_TO</type>
<position>106.5,-68</position>
<input>
<ID>IN_0</ID>682 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I2</lparam></gate>
<gate>
<ID>774</ID>
<type>DE_TO</type>
<position>108.5,-68</position>
<input>
<ID>IN_0</ID>683 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I3</lparam></gate>
<gate>
<ID>775</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>114,-61</position>
<input>
<ID>ENABLE_0</ID>693 </input>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>70 </input>
<output>
<ID>OUT_0</ID>684 </output>
<output>
<ID>OUT_1</ID>685 </output>
<output>
<ID>OUT_2</ID>686 </output>
<output>
<ID>OUT_3</ID>687 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>776</ID>
<type>DE_TO</type>
<position>111.5,-68</position>
<input>
<ID>IN_0</ID>684 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I4</lparam></gate>
<gate>
<ID>777</ID>
<type>DE_TO</type>
<position>113.5,-68</position>
<input>
<ID>IN_0</ID>685 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I5</lparam></gate>
<gate>
<ID>778</ID>
<type>DE_TO</type>
<position>115.5,-68</position>
<input>
<ID>IN_0</ID>686 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I6</lparam></gate>
<gate>
<ID>779</ID>
<type>DE_TO</type>
<position>117.5,-68</position>
<input>
<ID>IN_0</ID>687 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I7</lparam></gate>
<gate>
<ID>780</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>127.5,-61</position>
<input>
<ID>ENABLE_0</ID>700 </input>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>65 </input>
<input>
<ID>IN_3</ID>66 </input>
<output>
<ID>OUT_0</ID>688 </output>
<output>
<ID>OUT_1</ID>689 </output>
<output>
<ID>OUT_2</ID>690 </output>
<output>
<ID>OUT_3</ID>691 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>781</ID>
<type>DE_TO</type>
<position>125,-68</position>
<input>
<ID>IN_0</ID>688 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I8</lparam></gate>
<gate>
<ID>782</ID>
<type>DE_TO</type>
<position>127,-68</position>
<input>
<ID>IN_0</ID>689 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I9</lparam></gate>
<gate>
<ID>783</ID>
<type>DE_TO</type>
<position>129,-68</position>
<input>
<ID>IN_0</ID>690 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I10</lparam></gate>
<gate>
<ID>784</ID>
<type>DE_TO</type>
<position>131,-68</position>
<input>
<ID>IN_0</ID>691 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I11</lparam></gate>
<gate>
<ID>785</ID>
<type>DA_FROM</type>
<position>119,-61</position>
<input>
<ID>IN_0</ID>693 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID IR-PC</lparam></gate>
<gate>
<ID>786</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>138.5,-68</position>
<input>
<ID>ENABLE_0</ID>699 </input>
<input>
<ID>IN_0</ID>698 </input>
<input>
<ID>IN_1</ID>698 </input>
<input>
<ID>IN_2</ID>698 </input>
<input>
<ID>IN_3</ID>698 </input>
<output>
<ID>OUT_0</ID>694 </output>
<output>
<ID>OUT_1</ID>695 </output>
<output>
<ID>OUT_2</ID>696 </output>
<output>
<ID>OUT_3</ID>697 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>787</ID>
<type>DE_TO</type>
<position>136,-75</position>
<input>
<ID>IN_0</ID>694 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I8</lparam></gate>
<gate>
<ID>788</ID>
<type>DE_TO</type>
<position>138,-75</position>
<input>
<ID>IN_0</ID>695 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I9</lparam></gate>
<gate>
<ID>789</ID>
<type>DE_TO</type>
<position>140,-75</position>
<input>
<ID>IN_0</ID>696 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I10</lparam></gate>
<gate>
<ID>790</ID>
<type>DE_TO</type>
<position>142,-75</position>
<input>
<ID>IN_0</ID>697 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I11</lparam></gate>
<gate>
<ID>792</ID>
<type>BA_TRI_STATE</type>
<position>140,-63</position>
<input>
<ID>ENABLE_0</ID>699 </input>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>698 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>793</ID>
<type>DA_FROM</type>
<position>145.5,-68</position>
<input>
<ID>IN_0</ID>699 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PC EXS</lparam></gate>
<gate>
<ID>794</ID>
<type>DA_FROM</type>
<position>132.5,-59</position>
<input>
<ID>IN_0</ID>700 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCDIR</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>78,0.5</position>
<gparam>LABEL_TEXT Instruction Register and Decode stage 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>DE_TO</type>
<position>145,-31.5</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BNZ</lparam></gate>
<gate>
<ID>63</ID>
<type>AM_REGISTER16</type>
<position>33,-50</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>56 </input>
<input>
<ID>IN_10</ID>46 </input>
<input>
<ID>IN_11</ID>44 </input>
<input>
<ID>IN_12</ID>43 </input>
<input>
<ID>IN_13</ID>42 </input>
<input>
<ID>IN_14</ID>41 </input>
<input>
<ID>IN_15</ID>40 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>54 </input>
<input>
<ID>IN_4</ID>52 </input>
<input>
<ID>IN_5</ID>51 </input>
<input>
<ID>IN_6</ID>50 </input>
<input>
<ID>IN_7</ID>49 </input>
<input>
<ID>IN_8</ID>48 </input>
<input>
<ID>IN_9</ID>47 </input>
<output>
<ID>OUT_0</ID>71 </output>
<output>
<ID>OUT_1</ID>72 </output>
<output>
<ID>OUT_10</ID>65 </output>
<output>
<ID>OUT_11</ID>66 </output>
<output>
<ID>OUT_12</ID>59 </output>
<output>
<ID>OUT_13</ID>60 </output>
<output>
<ID>OUT_14</ID>61 </output>
<output>
<ID>OUT_15</ID>58 </output>
<output>
<ID>OUT_2</ID>73 </output>
<output>
<ID>OUT_3</ID>74 </output>
<output>
<ID>OUT_4</ID>67 </output>
<output>
<ID>OUT_5</ID>68 </output>
<output>
<ID>OUT_6</ID>69 </output>
<output>
<ID>OUT_7</ID>70 </output>
<output>
<ID>OUT_8</ID>63 </output>
<output>
<ID>OUT_9</ID>64 </output>
<input>
<ID>clear</ID>37 </input>
<input>
<ID>clock</ID>36 </input>
<input>
<ID>count_enable</ID>38 </input>
<input>
<ID>count_up</ID>38 </input>
<input>
<ID>load</ID>39 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 53539</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>34.5,-63.5</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>66</ID>
<type>FF_GND</type>
<position>34,-60.5</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>FF_GND</type>
<position>34,-38.5</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>70</ID>
<type>DA_FROM</type>
<position>32,-36</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>9.5,-21</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>10,-23.5</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>9.5,-27</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>76</ID>
<type>DA_FROM</type>
<position>10,-29.5</position>
<input>
<ID>IN_0</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>10,-32.5</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>11,-35</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>79</ID>
<type>DA_FROM</type>
<position>10,-38.5</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>10.5,-41</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>81</ID>
<type>DA_FROM</type>
<position>11.5,-45</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>12,-47.5</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>11,-50.5</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>12,-53.5</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>85</ID>
<type>DA_FROM</type>
<position>12,-55.5</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>664</ID>
<type>AE_DFF_LOW</type>
<position>5,-7.5</position>
<input>
<ID>IN_0</ID>584 </input>
<output>
<ID>OUTINV_0</ID>584 </output>
<output>
<ID>OUT_0</ID>587 </output>
<input>
<ID>clear</ID>583 </input>
<input>
<ID>clock</ID>586 </input>
<input>
<ID>set</ID>585 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>86</ID>
<type>DA_FROM</type>
<position>12,-58.5</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>87</ID>
<type>DA_FROM</type>
<position>11.5,-61.5</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>666</ID>
<type>EE_VDD</type>
<position>5,-2</position>
<output>
<ID>OUT_0</ID>585 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>88</ID>
<type>DA_FROM</type>
<position>11.5,-65.5</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>668</ID>
<type>EE_VDD</type>
<position>5,-13</position>
<output>
<ID>OUT_0</ID>583 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>90</ID>
<type>BI_DECODER_4x16</type>
<position>57.5,-26.5</position>
<input>
<ID>ENABLE</ID>62 </input>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>60 </input>
<input>
<ID>IN_2</ID>61 </input>
<input>
<ID>IN_3</ID>58 </input>
<output>
<ID>OUT_10</ID>1063 </output>
<output>
<ID>OUT_11</ID>1062 </output>
<output>
<ID>OUT_12</ID>579 </output>
<output>
<ID>OUT_13</ID>368 </output>
<output>
<ID>OUT_14</ID>261 </output>
<output>
<ID>OUT_15</ID>75 </output>
<output>
<ID>OUT_9</ID>1064 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>669</ID>
<type>DA_FROM</type>
<position>-3.5,-8.5</position>
<input>
<ID>IN_0</ID>586 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>92</ID>
<type>DA_FROM</type>
<position>46.5,-19</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Execute</lparam></gate>
<gate>
<ID>671</ID>
<type>DE_TO</type>
<position>15.5,-8.5</position>
<input>
<ID>IN_0</ID>584 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Execute</lparam></gate>
<gate>
<ID>93</ID>
<type>DE_TO</type>
<position>73.5,-83</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>94</ID>
<type>DE_TO</type>
<position>69.5,-83.5</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>673</ID>
<type>DE_TO</type>
<position>16.5,-5.5</position>
<input>
<ID>IN_0</ID>587 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>95</ID>
<type>DE_TO</type>
<position>66,-84</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>96</ID>
<type>DE_TO</type>
<position>63,-84</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>483</ID>
<type>DE_TO</type>
<position>94.5,-22</position>
<input>
<ID>IN_0</ID>579 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MOVEI</lparam></gate>
<gate>
<ID>97</ID>
<type>DE_TO</type>
<position>59.5,-84</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>291</ID>
<type>DE_TO</type>
<position>78,-20</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID JMP</lparam></gate>
<gate>
<ID>98</ID>
<type>DE_TO</type>
<position>56,-84</position>
<input>
<ID>IN_0</ID>110 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>99</ID>
<type>DE_TO</type>
<position>53,-84.5</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>293</ID>
<type>DE_TO</type>
<position>142,-28</position>
<input>
<ID>IN_0</ID>262 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZ</lparam></gate>
<gate>
<ID>100</ID>
<type>DE_TO</type>
<position>49.5,-84.5</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>101</ID>
<type>DE_TO</type>
<position>25,-85</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>102</ID>
<type>DE_TO</type>
<position>28.5,-85</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>31.5,-85</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>1069</ID>
<type>DE_TO</type>
<position>103,-23.5</position>
<input>
<ID>IN_0</ID>1062 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MOVE</lparam></gate>
<gate>
<ID>104</ID>
<type>DE_TO</type>
<position>34.5,-85</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>1070</ID>
<type>DE_TO</type>
<position>117.5,-24.5</position>
<input>
<ID>IN_0</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STORE</lparam></gate>
<gate>
<ID>105</ID>
<type>DE_TO</type>
<position>37.5,-85</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>1071</ID>
<type>DE_TO</type>
<position>107,-26.5</position>
<input>
<ID>IN_0</ID>1064 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>40,-85</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>1072</ID>
<type>DE_TO</type>
<position>169,-36.5</position>
<input>
<ID>IN_0</ID>1065 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STA</lparam></gate>
<gate>
<ID>107</ID>
<type>DE_TO</type>
<position>42.5,-84.5</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>1073</ID>
<type>DE_TO</type>
<position>167,-42.5</position>
<input>
<ID>IN_0</ID>1066 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STA+</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>46,-84.5</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>110</ID>
<type>BI_DECODER_4x16</type>
<position>135.5,-42</position>
<input>
<ID>ENABLE</ID>75 </input>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>65 </input>
<input>
<ID>IN_3</ID>66 </input>
<output>
<ID>OUT_13</ID>185 </output>
<output>
<ID>OUT_14</ID>262 </output>
<output>
<ID>OUT_15</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>112</ID>
<type>BI_DECODER_4x16</type>
<position>144,-46</position>
<input>
<ID>ENABLE</ID>76 </input>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>70 </input>
<output>
<ID>OUT_15</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>114</ID>
<type>BI_DECODER_4x16</type>
<position>158.5,-50</position>
<input>
<ID>ENABLE</ID>77 </input>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<output>
<ID>OUT_14</ID>1066 </output>
<output>
<ID>OUT_15</ID>1065 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>116</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>47,-73.5</position>
<input>
<ID>ENABLE_0</ID>125 </input>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_10</ID>65 </input>
<input>
<ID>IN_11</ID>66 </input>
<input>
<ID>IN_12</ID>111 </input>
<input>
<ID>IN_13</ID>111 </input>
<input>
<ID>IN_14</ID>111 </input>
<input>
<ID>IN_15</ID>111 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<input>
<ID>IN_4</ID>67 </input>
<input>
<ID>IN_5</ID>68 </input>
<input>
<ID>IN_6</ID>69 </input>
<input>
<ID>IN_7</ID>70 </input>
<input>
<ID>IN_8</ID>63 </input>
<input>
<ID>IN_9</ID>64 </input>
<output>
<ID>OUT_0</ID>99 </output>
<output>
<ID>OUT_1</ID>100 </output>
<output>
<ID>OUT_10</ID>110 </output>
<output>
<ID>OUT_11</ID>109 </output>
<output>
<ID>OUT_12</ID>98 </output>
<output>
<ID>OUT_13</ID>97 </output>
<output>
<ID>OUT_14</ID>96 </output>
<output>
<ID>OUT_15</ID>95 </output>
<output>
<ID>OUT_2</ID>101 </output>
<output>
<ID>OUT_3</ID>102 </output>
<output>
<ID>OUT_4</ID>103 </output>
<output>
<ID>OUT_5</ID>104 </output>
<output>
<ID>OUT_6</ID>105 </output>
<output>
<ID>OUT_7</ID>106 </output>
<output>
<ID>OUT_8</ID>107 </output>
<output>
<ID>OUT_9</ID>108 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>120</ID>
<type>BA_TRI_STATE</type>
<position>54.5,-67.5</position>
<input>
<ID>ENABLE_0</ID>94 </input>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>111 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>122</ID>
<type>EE_VDD</type>
<position>57.5,-65.5</position>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>126</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>67.5,-60.5</position>
<input>
<ID>ENABLE_0</ID>124 </input>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<output>
<ID>OUT_0</ID>112 </output>
<output>
<ID>OUT_1</ID>113 </output>
<output>
<ID>OUT_2</ID>114 </output>
<output>
<ID>OUT_3</ID>115 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>128</ID>
<type>DE_TO</type>
<position>65,-67.5</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 0</lparam></gate>
<gate>
<ID>129</ID>
<type>DE_TO</type>
<position>67,-67.5</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 1</lparam></gate>
<gate>
<ID>130</ID>
<type>DE_TO</type>
<position>69,-67.5</position>
<input>
<ID>IN_0</ID>114 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 2</lparam></gate>
<gate>
<ID>131</ID>
<type>DE_TO</type>
<position>71,-67.5</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 3</lparam></gate>
<gate>
<ID>132</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>76.5,-60.5</position>
<input>
<ID>ENABLE_0</ID>124 </input>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>70 </input>
<output>
<ID>OUT_0</ID>116 </output>
<output>
<ID>OUT_1</ID>117 </output>
<output>
<ID>OUT_2</ID>118 </output>
<output>
<ID>OUT_3</ID>119 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>133</ID>
<type>DE_TO</type>
<position>74,-67.5</position>
<input>
<ID>IN_0</ID>116 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 4</lparam></gate>
<gate>
<ID>134</ID>
<type>DE_TO</type>
<position>76,-67.5</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 5</lparam></gate>
<gate>
<ID>135</ID>
<type>DE_TO</type>
<position>78,-67.5</position>
<input>
<ID>IN_0</ID>118 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 6</lparam></gate>
<gate>
<ID>136</ID>
<type>DE_TO</type>
<position>80,-67.5</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 7</lparam></gate>
<gate>
<ID>137</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>86,-60.5</position>
<input>
<ID>ENABLE_0</ID>124 </input>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>65 </input>
<input>
<ID>IN_3</ID>66 </input>
<output>
<ID>OUT_0</ID>120 </output>
<output>
<ID>OUT_1</ID>121 </output>
<output>
<ID>OUT_2</ID>122 </output>
<output>
<ID>OUT_3</ID>123 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>138</ID>
<type>DE_TO</type>
<position>83.5,-67.5</position>
<input>
<ID>IN_0</ID>120 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 8</lparam></gate>
<gate>
<ID>139</ID>
<type>DE_TO</type>
<position>85.5,-67.5</position>
<input>
<ID>IN_0</ID>121 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 9</lparam></gate>
<gate>
<ID>140</ID>
<type>DE_TO</type>
<position>87.5,-67.5</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 10</lparam></gate>
<gate>
<ID>141</ID>
<type>DE_TO</type>
<position>89.5,-67.5</position>
<input>
<ID>IN_0</ID>123 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 11</lparam></gate>
<gate>
<ID>143</ID>
<type>DA_FROM</type>
<position>92.5,-60.5</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID IR-AD</lparam></gate>
<gate>
<ID>145</ID>
<type>DA_FROM</type>
<position>58.5,-73.5</position>
<input>
<ID>IN_0</ID>125 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Imm</lparam></gate>
<gate>
<ID>146</ID>
<type>DE_TO</type>
<position>114.5,-87</position>
<input>
<ID>IN_0</ID>126 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Ck2</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_TOGGLE</type>
<position>123.5,-87</position>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>378</ID>
<type>DE_TO</type>
<position>86.5,-21</position>
<input>
<ID>IN_0</ID>368 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADDI</lparam></gate>
<gate>
<ID>770</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>105,-61</position>
<input>
<ID>ENABLE_0</ID>693 </input>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<output>
<ID>OUT_0</ID>680 </output>
<output>
<ID>OUT_1</ID>681 </output>
<output>
<ID>OUT_2</ID>682 </output>
<output>
<ID>OUT_3</ID>683 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>771</ID>
<type>DE_TO</type>
<position>102.5,-68</position>
<input>
<ID>IN_0</ID>680 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I0</lparam></gate>
<wire>
<ID>579</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-22,92.5,-22</points>
<connection>
<GID>90</GID>
<name>OUT_12</name></connection>
<connection>
<GID>483</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-12,5,-11.5</points>
<connection>
<GID>664</GID>
<name>clear</name></connection>
<connection>
<GID>668</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-8.5,11,2.5</points>
<intersection>-8.5 2</intersection>
<intersection>2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,2.5,11,2.5</points>
<intersection>2 3</intersection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-8.5,13.5,-8.5</points>
<connection>
<GID>664</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>2,-5.5,2,2.5</points>
<connection>
<GID>664</GID>
<name>IN_0</name></connection>
<intersection>2.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-3.5,5,-3</points>
<connection>
<GID>666</GID>
<name>OUT_0</name></connection>
<connection>
<GID>664</GID>
<name>set</name></connection></vsegment></shape></wire>
<wire>
<ID>586</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-8.5,2,-8.5</points>
<connection>
<GID>664</GID>
<name>clock</name></connection>
<connection>
<GID>669</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8,-5.5,14.5,-5.5</points>
<connection>
<GID>664</GID>
<name>OUT_0</name></connection>
<connection>
<GID>673</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-63.5,32,-59.5</points>
<connection>
<GID>63</GID>
<name>clock</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-63.5,32.5,-63.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-59.5,34,-59.5</points>
<connection>
<GID>63</GID>
<name>clear</name></connection>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-40.5,34,-39.5</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>-40.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>33,-40.5,34,-40.5</points>
<connection>
<GID>63</GID>
<name>count_up</name></connection>
<connection>
<GID>63</GID>
<name>count_enable</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-40.5,32,-38</points>
<connection>
<GID>63</GID>
<name>load</name></connection>
<connection>
<GID>70</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-21,27.5,-21</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>27.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27.5,-42.5,27.5,-21</points>
<intersection>-42.5 4</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>27.5,-42.5,28,-42.5</points>
<connection>
<GID>63</GID>
<name>IN_15</name></connection>
<intersection>27.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-43.5,26,-23.5</points>
<intersection>-43.5 1</intersection>
<intersection>-23.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-43.5,28,-43.5</points>
<connection>
<GID>63</GID>
<name>IN_14</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>12,-23.5,26,-23.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-44.5,24,-27</points>
<intersection>-44.5 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-44.5,28,-44.5</points>
<connection>
<GID>63</GID>
<name>IN_13</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-27,24,-27</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-45.5,22,-29.5</points>
<intersection>-45.5 1</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-45.5,28,-45.5</points>
<connection>
<GID>63</GID>
<name>IN_12</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-29.5,22,-29.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-46.5,21,-32.5</points>
<intersection>-46.5 1</intersection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-46.5,28,-46.5</points>
<connection>
<GID>63</GID>
<name>IN_11</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-32.5,21,-32.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-47.5,20.5,-35</points>
<intersection>-47.5 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-47.5,28,-47.5</points>
<connection>
<GID>63</GID>
<name>IN_10</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-35,20.5,-35</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-48.5,20,-38.5</points>
<intersection>-48.5 1</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-48.5,28,-48.5</points>
<connection>
<GID>63</GID>
<name>IN_9</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-38.5,20,-38.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-49.5,20,-41</points>
<intersection>-49.5 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-49.5,28,-49.5</points>
<connection>
<GID>63</GID>
<name>IN_8</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-41,20,-41</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-50.5,19.5,-45</points>
<intersection>-50.5 1</intersection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-50.5,28,-50.5</points>
<connection>
<GID>63</GID>
<name>IN_7</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-45,19.5,-45</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-51.5,18.5,-47.5</points>
<intersection>-51.5 1</intersection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-51.5,28,-51.5</points>
<connection>
<GID>63</GID>
<name>IN_6</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-47.5,18.5,-47.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-52.5,17.5,-50.5</points>
<intersection>-52.5 1</intersection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-52.5,28,-52.5</points>
<connection>
<GID>63</GID>
<name>IN_5</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-50.5,17.5,-50.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-53.5,28,-53.5</points>
<connection>
<GID>63</GID>
<name>IN_4</name></connection>
<connection>
<GID>84</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-55.5,23.5,-55.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>23.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>23.5,-55.5,23.5,-54.5</points>
<intersection>-55.5 1</intersection>
<intersection>-54.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>23.5,-54.5,28,-54.5</points>
<connection>
<GID>63</GID>
<name>IN_3</name></connection>
<intersection>23.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-58.5,25,-55.5</points>
<intersection>-58.5 2</intersection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-55.5,28,-55.5</points>
<connection>
<GID>63</GID>
<name>IN_2</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-58.5,25,-58.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-61.5,26,-56.5</points>
<intersection>-61.5 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-56.5,28,-56.5</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-61.5,26,-61.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-65.5,27.5,-57.5</points>
<intersection>-65.5 2</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-57.5,28,-57.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-65.5,27.5,-65.5</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-31,54.5,-31</points>
<connection>
<GID>90</GID>
<name>IN_3</name></connection>
<intersection>48 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>48,-42.5,48,-31</points>
<intersection>-42.5 5</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38,-42.5,48,-42.5</points>
<connection>
<GID>63</GID>
<name>OUT_15</name></connection>
<intersection>48 4</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-34,54.5,-34</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>53.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>53.5,-45.5,53.5,-34</points>
<intersection>-45.5 5</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38,-45.5,53.5,-45.5</points>
<connection>
<GID>63</GID>
<name>OUT_12</name></connection>
<intersection>53.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-33,54.5,-33</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<intersection>51.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-44.5,51.5,-33</points>
<intersection>-44.5 5</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38,-44.5,51.5,-44.5</points>
<connection>
<GID>63</GID>
<name>OUT_13</name></connection>
<intersection>51.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-32,54.5,-32</points>
<connection>
<GID>90</GID>
<name>IN_2</name></connection>
<intersection>50 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>50,-43.5,50,-32</points>
<intersection>-43.5 5</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38,-43.5,50,-43.5</points>
<connection>
<GID>63</GID>
<name>OUT_14</name></connection>
<intersection>50 4</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-19,54.5,-19</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<connection>
<GID>90</GID>
<name>ENABLE</name></connection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-49.5,132.5,-49.5</points>
<connection>
<GID>63</GID>
<name>OUT_8</name></connection>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>47.5 13</intersection>
<intersection>84.5 16</intersection>
<intersection>126 20</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>47.5,-71.5,47.5,-49.5</points>
<connection>
<GID>116</GID>
<name>IN_8</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>84.5,-58.5,84.5,-49.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>126,-59,126,-49.5</points>
<connection>
<GID>780</GID>
<name>IN_0</name></connection>
<intersection>-49.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-48.5,132.5,-48.5</points>
<connection>
<GID>63</GID>
<name>OUT_9</name></connection>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>48.5 13</intersection>
<intersection>85.5 23</intersection>
<intersection>127 27</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>48.5,-71.5,48.5,-48.5</points>
<connection>
<GID>116</GID>
<name>IN_9</name></connection>
<intersection>-48.5 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>85.5,-58.5,85.5,-48.5</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<intersection>-48.5 1</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>127,-59,127,-48.5</points>
<connection>
<GID>780</GID>
<name>IN_1</name></connection>
<intersection>-48.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-47.5,132.5,-47.5</points>
<connection>
<GID>63</GID>
<name>OUT_10</name></connection>
<connection>
<GID>110</GID>
<name>IN_2</name></connection>
<intersection>49.5 13</intersection>
<intersection>86.5 22</intersection>
<intersection>128 26</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>49.5,-71.5,49.5,-47.5</points>
<connection>
<GID>116</GID>
<name>IN_10</name></connection>
<intersection>-47.5 1</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>86.5,-58.5,86.5,-47.5</points>
<connection>
<GID>137</GID>
<name>IN_2</name></connection>
<intersection>-47.5 1</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>128,-59,128,-47.5</points>
<connection>
<GID>780</GID>
<name>IN_2</name></connection>
<intersection>-47.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-46.5,132.5,-46.5</points>
<connection>
<GID>63</GID>
<name>OUT_11</name></connection>
<connection>
<GID>110</GID>
<name>IN_3</name></connection>
<intersection>50.5 13</intersection>
<intersection>87.5 27</intersection>
<intersection>129 31</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>50.5,-71.5,50.5,-46.5</points>
<connection>
<GID>116</GID>
<name>IN_11</name></connection>
<intersection>-64.5 15</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>50.5,-64.5,54.5,-64.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>50.5 13</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>87.5,-58.5,87.5,-46.5</points>
<connection>
<GID>137</GID>
<name>IN_3</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>129,-59,129,-46.5</points>
<connection>
<GID>780</GID>
<name>IN_3</name></connection>
<intersection>-46.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-53.5,141,-53.5</points>
<connection>
<GID>63</GID>
<name>OUT_4</name></connection>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>43.5 4</intersection>
<intersection>75 8</intersection>
<intersection>112.5 15</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>43.5,-71.5,43.5,-53.5</points>
<connection>
<GID>116</GID>
<name>IN_4</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>75,-58.5,75,-53.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>112.5,-59,112.5,-53.5</points>
<connection>
<GID>775</GID>
<name>IN_0</name></connection>
<intersection>-53.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-20,76,-20</points>
<connection>
<GID>90</GID>
<name>OUT_14</name></connection>
<connection>
<GID>291</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-52.5,141,-52.5</points>
<connection>
<GID>63</GID>
<name>OUT_5</name></connection>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>44.5 4</intersection>
<intersection>76 8</intersection>
<intersection>113.5 15</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>44.5,-71.5,44.5,-52.5</points>
<connection>
<GID>116</GID>
<name>IN_5</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>76,-58.5,76,-52.5</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>113.5,-59,113.5,-52.5</points>
<connection>
<GID>775</GID>
<name>IN_1</name></connection>
<intersection>-52.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-35.5,139,-28</points>
<intersection>-35.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,-35.5,139,-35.5</points>
<connection>
<GID>110</GID>
<name>OUT_14</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139,-28,140,-28</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-51.5,141,-51.5</points>
<connection>
<GID>63</GID>
<name>OUT_6</name></connection>
<connection>
<GID>112</GID>
<name>IN_2</name></connection>
<intersection>45.5 4</intersection>
<intersection>77 8</intersection>
<intersection>114.5 15</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>45.5,-71.5,45.5,-51.5</points>
<connection>
<GID>116</GID>
<name>IN_6</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>77,-58.5,77,-51.5</points>
<connection>
<GID>132</GID>
<name>IN_2</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>114.5,-59,114.5,-51.5</points>
<connection>
<GID>775</GID>
<name>IN_2</name></connection>
<intersection>-51.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-50.5,141,-50.5</points>
<connection>
<GID>63</GID>
<name>OUT_7</name></connection>
<connection>
<GID>112</GID>
<name>IN_3</name></connection>
<intersection>46.5 4</intersection>
<intersection>78 8</intersection>
<intersection>115.5 15</intersection>
<intersection>140 16</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>46.5,-71.5,46.5,-50.5</points>
<connection>
<GID>116</GID>
<name>IN_7</name></connection>
<intersection>-50.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>78,-58.5,78,-50.5</points>
<connection>
<GID>132</GID>
<name>IN_3</name></connection>
<intersection>-50.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>115.5,-59,115.5,-50.5</points>
<connection>
<GID>775</GID>
<name>IN_3</name></connection>
<intersection>-50.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>140,-60,140,-50.5</points>
<connection>
<GID>792</GID>
<name>IN_0</name></connection>
<intersection>-50.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-57.5,155.5,-57.5</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>39.5 7</intersection>
<intersection>66 8</intersection>
<intersection>103.5 12</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>39.5,-71.5,39.5,-57.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>-57.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>66,-58.5,66,-57.5</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-57.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>103.5,-59,103.5,-57.5</points>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<intersection>-57.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-56.5,155.5,-56.5</points>
<connection>
<GID>63</GID>
<name>OUT_1</name></connection>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>40.5 7</intersection>
<intersection>67 9</intersection>
<intersection>104.5 13</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>40.5,-71.5,40.5,-56.5</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>67,-58.5,67,-56.5</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>104.5,-59,104.5,-56.5</points>
<connection>
<GID>770</GID>
<name>IN_1</name></connection>
<intersection>-56.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-55.5,155.5,-55.5</points>
<connection>
<GID>63</GID>
<name>OUT_2</name></connection>
<connection>
<GID>114</GID>
<name>IN_2</name></connection>
<intersection>41.5 7</intersection>
<intersection>68 8</intersection>
<intersection>105.5 12</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>41.5,-71.5,41.5,-55.5</points>
<connection>
<GID>116</GID>
<name>IN_2</name></connection>
<intersection>-55.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>68,-58.5,68,-55.5</points>
<connection>
<GID>126</GID>
<name>IN_2</name></connection>
<intersection>-55.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>105.5,-59,105.5,-55.5</points>
<connection>
<GID>770</GID>
<name>IN_2</name></connection>
<intersection>-55.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-54.5,155.5,-54.5</points>
<connection>
<GID>63</GID>
<name>OUT_3</name></connection>
<connection>
<GID>114</GID>
<name>IN_3</name></connection>
<intersection>42.5 7</intersection>
<intersection>69 8</intersection>
<intersection>106.5 12</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>42.5,-71.5,42.5,-54.5</points>
<connection>
<GID>116</GID>
<name>IN_3</name></connection>
<intersection>-54.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>69,-58.5,69,-54.5</points>
<connection>
<GID>126</GID>
<name>IN_3</name></connection>
<intersection>-54.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>106.5,-59,106.5,-54.5</points>
<connection>
<GID>770</GID>
<name>IN_3</name></connection>
<intersection>-54.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-34.5,73.5,-19</points>
<intersection>-34.5 5</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>60.5,-19,73.5,-19</points>
<connection>
<GID>90</GID>
<name>OUT_15</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>73.5,-34.5,132.5,-34.5</points>
<connection>
<GID>110</GID>
<name>ENABLE</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-38.5,140,-34.5</points>
<intersection>-38.5 3</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>138.5,-34.5,140,-34.5</points>
<connection>
<GID>110</GID>
<name>OUT_15</name></connection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>140,-38.5,141,-38.5</points>
<connection>
<GID>112</GID>
<name>ENABLE</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150.5,-42.5,150.5,-38.5</points>
<intersection>-42.5 1</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-42.5,155.5,-42.5</points>
<connection>
<GID>114</GID>
<name>ENABLE</name></connection>
<intersection>150.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147,-38.5,150.5,-38.5</points>
<connection>
<GID>112</GID>
<name>OUT_15</name></connection>
<intersection>150.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-67.5,57.5,-66.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-67.5,57.5,-67.5</points>
<connection>
<GID>120</GID>
<name>ENABLE_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-81,73.5,-75.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>-75.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-75.5,73.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_15</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-81.5,69.5,-76.5</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>-76.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>53.5,-76.5,53.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_14</name></connection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-76.5,69.5,-76.5</points>
<intersection>53.5 1</intersection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-82,66,-77.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>-77.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>52.5,-77.5,52.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_13</name></connection>
<intersection>-77.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>52.5,-77.5,66,-77.5</points>
<intersection>52.5 1</intersection>
<intersection>66 0</intersection></hsegment></shape></wire>
<wire>
<ID>1062</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-23.5,80.5,-23</points>
<intersection>-23.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-23,80.5,-23</points>
<connection>
<GID>90</GID>
<name>OUT_11</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80.5,-23.5,101,-23.5</points>
<connection>
<GID>1069</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-82,63,-78</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>-78 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>51.5,-78,51.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_12</name></connection>
<intersection>-78 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-78,63,-78</points>
<intersection>51.5 1</intersection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>1063</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-24.5,79.5,-24</points>
<intersection>-24.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-24,79.5,-24</points>
<connection>
<GID>90</GID>
<name>OUT_10</name></connection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79.5,-24.5,115.5,-24.5</points>
<connection>
<GID>1070</GID>
<name>IN_0</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>25,-83,25,-76</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-76 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25,-76,39.5,-76</points>
<intersection>25 1</intersection>
<intersection>39.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>39.5,-76,39.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<intersection>-76 2</intersection></vsegment></shape></wire>
<wire>
<ID>1064</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-26.5,82.5,-25</points>
<intersection>-26.5 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-25,82.5,-25</points>
<connection>
<GID>90</GID>
<name>OUT_9</name></connection>
<intersection>82.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-26.5,105,-26.5</points>
<connection>
<GID>1071</GID>
<name>IN_0</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1065</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161.5,-36.5,167,-36.5</points>
<connection>
<GID>1072</GID>
<name>IN_0</name></connection>
<intersection>161.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>161.5,-42.5,161.5,-36.5</points>
<connection>
<GID>114</GID>
<name>OUT_15</name></connection>
<intersection>-36.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-83,28.5,-77</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>-77 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>40.5,-77,40.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_1</name></connection>
<intersection>-77 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-77,40.5,-77</points>
<intersection>28.5 0</intersection>
<intersection>40.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>680</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-66,102.5,-63</points>
<connection>
<GID>771</GID>
<name>IN_0</name></connection>
<intersection>-63 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>102.5,-63,103.5,-63</points>
<connection>
<GID>770</GID>
<name>OUT_0</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1066</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-43.5,163,-42.5</points>
<intersection>-43.5 1</intersection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161.5,-43.5,163,-43.5</points>
<connection>
<GID>114</GID>
<name>OUT_14</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163,-42.5,165,-42.5</points>
<connection>
<GID>1073</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-83,31.5,-78</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>-78 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>41.5,-78,41.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_2</name></connection>
<intersection>-78 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-78,41.5,-78</points>
<intersection>31.5 0</intersection>
<intersection>41.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-83,34.5,-78.5</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>-78.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>42.5,-78.5,42.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_3</name></connection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-78.5,42.5,-78.5</points>
<intersection>34.5 0</intersection>
<intersection>42.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>681</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-66,104.5,-63</points>
<connection>
<GID>770</GID>
<name>OUT_1</name></connection>
<connection>
<GID>772</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-83,37.5,-79</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>-79 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>43.5,-79,43.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_4</name></connection>
<intersection>-79 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-79,43.5,-79</points>
<intersection>37.5 0</intersection>
<intersection>43.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>682</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-66,105.5,-63</points>
<connection>
<GID>770</GID>
<name>OUT_2</name></connection>
<intersection>-66 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>105.5,-66,106.5,-66</points>
<connection>
<GID>773</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-83,40,-79.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>-79.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>44.5,-79.5,44.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_5</name></connection>
<intersection>-79.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>40,-79.5,44.5,-79.5</points>
<intersection>40 0</intersection>
<intersection>44.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>683</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-63.5,106.5,-63</points>
<connection>
<GID>770</GID>
<name>OUT_3</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>108.5,-66,108.5,-63.5</points>
<connection>
<GID>774</GID>
<name>IN_0</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>106.5,-63.5,108.5,-63.5</points>
<intersection>106.5 0</intersection>
<intersection>108.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-82.5,42.5,-80</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>-80 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>45.5,-80,45.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_6</name></connection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-80,45.5,-80</points>
<intersection>42.5 0</intersection>
<intersection>45.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>684</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-66,111.5,-63</points>
<connection>
<GID>776</GID>
<name>IN_0</name></connection>
<intersection>-63 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>111.5,-63,112.5,-63</points>
<connection>
<GID>775</GID>
<name>OUT_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-82.5,46,-79</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-79 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>46.5,-79,46.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_7</name></connection>
<intersection>-79 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>46,-79,46.5,-79</points>
<intersection>46 0</intersection>
<intersection>46.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>685</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-66,113.5,-63</points>
<connection>
<GID>777</GID>
<name>IN_0</name></connection>
<connection>
<GID>775</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-82.5,49.5,-81</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>-81 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>47.5,-81,47.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_8</name></connection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47.5,-81,49.5,-81</points>
<intersection>47.5 1</intersection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>686</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-66,115.5,-64.5</points>
<connection>
<GID>778</GID>
<name>IN_0</name></connection>
<intersection>-64.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>114.5,-64.5,115.5,-64.5</points>
<intersection>114.5 5</intersection>
<intersection>115.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>114.5,-64.5,114.5,-63</points>
<connection>
<GID>775</GID>
<name>OUT_2</name></connection>
<intersection>-64.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-82.5,53,-80</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>-80 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>48.5,-80,48.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_9</name></connection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-80,53,-80</points>
<intersection>48.5 1</intersection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>687</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>117.5,-66,117.5,-63</points>
<connection>
<GID>779</GID>
<name>IN_0</name></connection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115.5,-63,117.5,-63</points>
<connection>
<GID>775</GID>
<name>OUT_3</name></connection>
<intersection>117.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-82,59.5,-78.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>-78.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>50.5,-78.5,50.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_11</name></connection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-78.5,59.5,-78.5</points>
<intersection>50.5 1</intersection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>688</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-66,125,-63</points>
<connection>
<GID>781</GID>
<name>IN_0</name></connection>
<intersection>-63 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>125,-63,126,-63</points>
<connection>
<GID>780</GID>
<name>OUT_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-82,56,-79</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>-79 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>49.5,-79,49.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_10</name></connection>
<intersection>-79 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-79,56,-79</points>
<intersection>49.5 1</intersection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-66,127,-63</points>
<connection>
<GID>782</GID>
<name>IN_0</name></connection>
<connection>
<GID>780</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-71.5,54.5,-70</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<connection>
<GID>116</GID>
<name>IN_15</name></connection>
<intersection>-71.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>51.5,-71.5,54.5,-71.5</points>
<connection>
<GID>116</GID>
<name>IN_14</name></connection>
<connection>
<GID>116</GID>
<name>IN_13</name></connection>
<connection>
<GID>116</GID>
<name>IN_12</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>690</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-66,128,-63</points>
<connection>
<GID>780</GID>
<name>OUT_2</name></connection>
<intersection>-66 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>128,-66,129,-66</points>
<connection>
<GID>783</GID>
<name>IN_0</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-65.5,65,-62.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-62.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>65,-62.5,66,-62.5</points>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-63.5,129,-63</points>
<connection>
<GID>780</GID>
<name>OUT_3</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>131,-66,131,-63.5</points>
<connection>
<GID>784</GID>
<name>IN_0</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>129,-63.5,131,-63.5</points>
<intersection>129 0</intersection>
<intersection>131 1</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-65.5,67,-62.5</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<connection>
<GID>126</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-65.5,69,-62.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-62.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>68,-62.5,69,-62.5</points>
<connection>
<GID>126</GID>
<name>OUT_2</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>693</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-61,117,-61</points>
<connection>
<GID>775</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>785</GID>
<name>IN_0</name></connection>
<connection>
<GID>770</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-63,69,-62.5</points>
<connection>
<GID>126</GID>
<name>OUT_3</name></connection>
<intersection>-63 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>71,-65.5,71,-63</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69,-63,71,-63</points>
<intersection>69 0</intersection>
<intersection>71 1</intersection></hsegment></shape></wire>
<wire>
<ID>694</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-73,136,-70</points>
<connection>
<GID>787</GID>
<name>IN_0</name></connection>
<intersection>-70 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>136,-70,137,-70</points>
<connection>
<GID>786</GID>
<name>OUT_0</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-65.5,74,-62.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>-62.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>74,-62.5,75,-62.5</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>695</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-73,138,-70</points>
<connection>
<GID>786</GID>
<name>OUT_1</name></connection>
<connection>
<GID>788</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-65.5,76,-62.5</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<connection>
<GID>132</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>696</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-73,139,-70</points>
<connection>
<GID>786</GID>
<name>OUT_2</name></connection>
<intersection>-73 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>139,-73,140,-73</points>
<connection>
<GID>789</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-65.5,78,-64</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>-64 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-64,78,-64</points>
<intersection>77 5</intersection>
<intersection>78 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>77,-64,77,-62.5</points>
<connection>
<GID>132</GID>
<name>OUT_2</name></connection>
<intersection>-64 3</intersection></vsegment></shape></wire>
<wire>
<ID>697</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-70.5,140,-70</points>
<connection>
<GID>786</GID>
<name>OUT_3</name></connection>
<intersection>-70.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>142,-73,142,-70.5</points>
<connection>
<GID>790</GID>
<name>IN_0</name></connection>
<intersection>-70.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>140,-70.5,142,-70.5</points>
<intersection>140 0</intersection>
<intersection>142 1</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>80,-65.5,80,-62.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>78,-62.5,80,-62.5</points>
<connection>
<GID>132</GID>
<name>OUT_3</name></connection>
<intersection>80 1</intersection></hsegment></shape></wire>
<wire>
<ID>698</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-66,140,-65.5</points>
<connection>
<GID>792</GID>
<name>OUT_0</name></connection>
<intersection>-66 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>137,-66,140,-66</points>
<connection>
<GID>786</GID>
<name>IN_3</name></connection>
<connection>
<GID>786</GID>
<name>IN_2</name></connection>
<connection>
<GID>786</GID>
<name>IN_1</name></connection>
<connection>
<GID>786</GID>
<name>IN_0</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-65.5,83.5,-62.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-62.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>83.5,-62.5,84.5,-62.5</points>
<connection>
<GID>137</GID>
<name>OUT_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>699</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-68,143.5,-68</points>
<connection>
<GID>786</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>793</GID>
<name>IN_0</name></connection>
<intersection>143.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>143.5,-68,143.5,-63</points>
<intersection>-68 1</intersection>
<intersection>-63 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>142,-63,143.5,-63</points>
<connection>
<GID>792</GID>
<name>ENABLE_0</name></connection>
<intersection>143.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-65.5,85.5,-62.5</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<connection>
<GID>137</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-61,130.5,-59</points>
<connection>
<GID>780</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>794</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-65.5,87.5,-62.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>-62.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>86.5,-62.5,87.5,-62.5</points>
<connection>
<GID>137</GID>
<name>OUT_2</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-63,87.5,-62.5</points>
<connection>
<GID>137</GID>
<name>OUT_3</name></connection>
<intersection>-63 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>89.5,-65.5,89.5,-63</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-63,89.5,-63</points>
<intersection>87.5 0</intersection>
<intersection>89.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-60.5,90.5,-60.5</points>
<connection>
<GID>137</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>126</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>132</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>143</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-73.5,56.5,-73.5</points>
<connection>
<GID>116</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>145</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116.5,-87,121.5,-87</points>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection>
<connection>
<GID>146</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-21,84.5,-21</points>
<connection>
<GID>90</GID>
<name>OUT_13</name></connection>
<connection>
<GID>378</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140.5,-36.5,140.5,-31.5</points>
<intersection>-36.5 1</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,-36.5,140.5,-36.5</points>
<connection>
<GID>110</GID>
<name>OUT_13</name></connection>
<intersection>140.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140.5,-31.5,143,-31.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>140.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-33.0077,34.0073,1061.21,-593.759</PageViewport>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>166.5,-56</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>160.5,-55</position>
<input>
<ID>IN_0</ID>366 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>414</ID>
<type>DE_OR8</type>
<position>132,-255.5</position>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_1</ID>452 </input>
<input>
<ID>IN_2</ID>453 </input>
<input>
<ID>IN_3</ID>454 </input>
<input>
<ID>IN_4</ID>504 </input>
<input>
<ID>IN_5</ID>503 </input>
<input>
<ID>IN_6</ID>502 </input>
<input>
<ID>IN_7</ID>501 </input>
<output>
<ID>OUT</ID>525 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>415</ID>
<type>DA_FROM</type>
<position>122,-248.5</position>
<input>
<ID>IN_0</ID>451 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MOVEI</lparam></gate>
<gate>
<ID>416</ID>
<type>DA_FROM</type>
<position>114,-251</position>
<input>
<ID>IN_0</ID>452 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MOVE</lparam></gate>
<gate>
<ID>417</ID>
<type>DA_FROM</type>
<position>112.5,-253.5</position>
<input>
<ID>IN_0</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>829</ID>
<type>AA_LABEL</type>
<position>365.5,-40.5</position>
<gparam>LABEL_TEXT Address Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>830</ID>
<type>DE_OR8</type>
<position>392.5,-128</position>
<input>
<ID>IN_0</ID>816 </input>
<input>
<ID>IN_1</ID>817 </input>
<input>
<ID>IN_2</ID>818 </input>
<input>
<ID>IN_3</ID>819 </input>
<input>
<ID>IN_4</ID>823 </input>
<input>
<ID>IN_5</ID>822 </input>
<input>
<ID>IN_6</ID>821 </input>
<input>
<ID>IN_7</ID>820 </input>
<output>
<ID>OUT</ID>824 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>831</ID>
<type>DA_FROM</type>
<position>382.5,-121</position>
<input>
<ID>IN_0</ID>816 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>832</ID>
<type>DA_FROM</type>
<position>374.5,-123.5</position>
<input>
<ID>IN_0</ID>817 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>833</ID>
<type>DA_FROM</type>
<position>373,-126</position>
<input>
<ID>IN_0</ID>818 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>444</ID>
<type>DA_FROM</type>
<position>112.5,-256</position>
<input>
<ID>IN_0</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>834</ID>
<type>DA_FROM</type>
<position>373,-128.5</position>
<input>
<ID>IN_0</ID>819 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>445</ID>
<type>DE_OR8</type>
<position>132,-221</position>
<input>
<ID>IN_0</ID>526 </input>
<input>
<ID>IN_1</ID>527 </input>
<input>
<ID>IN_2</ID>528 </input>
<input>
<ID>IN_3</ID>529 </input>
<input>
<ID>IN_4</ID>576 </input>
<input>
<ID>IN_5</ID>575 </input>
<input>
<ID>IN_6</ID>574 </input>
<input>
<ID>IN_7</ID>530 </input>
<output>
<ID>OUT</ID>577 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>56</ID>
<type>DA_FROM</type>
<position>153.5,-57</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BNZ</lparam></gate>
<gate>
<ID>835</ID>
<type>DA_FROM</type>
<position>373,-131.5</position>
<input>
<ID>IN_0</ID>820 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>446</ID>
<type>DA_FROM</type>
<position>112.5,-259</position>
<input>
<ID>IN_0</ID>501 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>836</ID>
<type>DA_FROM</type>
<position>373,-134</position>
<input>
<ID>IN_0</ID>821 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>447</ID>
<type>DA_FROM</type>
<position>122,-214</position>
<input>
<ID>IN_0</ID>526 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADDI</lparam></gate>
<gate>
<ID>837</ID>
<type>DA_FROM</type>
<position>373.5,-137</position>
<input>
<ID>IN_0</ID>822 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>448</ID>
<type>DA_FROM</type>
<position>112.5,-261.5</position>
<input>
<ID>IN_0</ID>502 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>838</ID>
<type>DA_FROM</type>
<position>373.5,-139.5</position>
<input>
<ID>IN_0</ID>823 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>449</ID>
<type>DA_FROM</type>
<position>114,-216.5</position>
<input>
<ID>IN_0</ID>527 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>839</ID>
<type>DE_TO</type>
<position>402,-128</position>
<input>
<ID>IN_0</ID>824 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BUS-ADREG</lparam></gate>
<gate>
<ID>840</ID>
<type>DE_OR8</type>
<position>390,-62</position>
<input>
<ID>IN_0</ID>825 </input>
<input>
<ID>IN_1</ID>826 </input>
<input>
<ID>IN_2</ID>827 </input>
<input>
<ID>IN_3</ID>828 </input>
<input>
<ID>IN_4</ID>832 </input>
<input>
<ID>IN_5</ID>831 </input>
<input>
<ID>IN_6</ID>830 </input>
<input>
<ID>IN_7</ID>829 </input>
<output>
<ID>OUT</ID>833 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>841</ID>
<type>DA_FROM</type>
<position>380,-55</position>
<input>
<ID>IN_0</ID>825 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STA+</lparam></gate>
<gate>
<ID>842</ID>
<type>DA_FROM</type>
<position>372,-57.5</position>
<input>
<ID>IN_0</ID>826 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>843</ID>
<type>DA_FROM</type>
<position>370.5,-60</position>
<input>
<ID>IN_0</ID>827 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>844</ID>
<type>DA_FROM</type>
<position>370.5,-62.5</position>
<input>
<ID>IN_0</ID>828 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>845</ID>
<type>DA_FROM</type>
<position>370.5,-65.5</position>
<input>
<ID>IN_0</ID>829 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>456</ID>
<type>DA_FROM</type>
<position>113,-264.5</position>
<input>
<ID>IN_0</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>846</ID>
<type>DA_FROM</type>
<position>370.5,-68</position>
<input>
<ID>IN_0</ID>830 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>457</ID>
<type>DA_FROM</type>
<position>112.5,-219</position>
<input>
<ID>IN_0</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>847</ID>
<type>DA_FROM</type>
<position>371,-71</position>
<input>
<ID>IN_0</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>458</ID>
<type>DA_FROM</type>
<position>113,-267</position>
<input>
<ID>IN_0</ID>504 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>848</ID>
<type>DA_FROM</type>
<position>371,-73.5</position>
<input>
<ID>IN_0</ID>832 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>459</ID>
<type>DA_FROM</type>
<position>112.5,-221.5</position>
<input>
<ID>IN_0</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>849</ID>
<type>DE_TO</type>
<position>399.5,-62</position>
<input>
<ID>IN_0</ID>833 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INC-ADREG</lparam></gate>
<gate>
<ID>460</ID>
<type>DE_TO</type>
<position>141.5,-255.5</position>
<input>
<ID>IN_0</ID>525 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus-Acc</lparam></gate>
<gate>
<ID>850</ID>
<type>DE_OR8</type>
<position>390,-93.5</position>
<input>
<ID>IN_0</ID>834 </input>
<input>
<ID>IN_1</ID>835 </input>
<input>
<ID>IN_2</ID>836 </input>
<input>
<ID>IN_3</ID>837 </input>
<input>
<ID>IN_4</ID>841 </input>
<input>
<ID>IN_5</ID>840 </input>
<input>
<ID>IN_6</ID>839 </input>
<input>
<ID>IN_7</ID>838 </input>
<output>
<ID>OUT</ID>842 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>461</ID>
<type>DA_FROM</type>
<position>112.5,-224.5</position>
<input>
<ID>IN_0</ID>530 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>851</ID>
<type>DA_FROM</type>
<position>380,-86.5</position>
<input>
<ID>IN_0</ID>834 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>852</ID>
<type>DA_FROM</type>
<position>372,-89</position>
<input>
<ID>IN_0</ID>835 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>463</ID>
<type>DA_FROM</type>
<position>112.5,-227</position>
<input>
<ID>IN_0</ID>574 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>853</ID>
<type>DA_FROM</type>
<position>370.5,-91.5</position>
<input>
<ID>IN_0</ID>836 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>854</ID>
<type>DA_FROM</type>
<position>370.5,-94</position>
<input>
<ID>IN_0</ID>837 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>855</ID>
<type>DA_FROM</type>
<position>370.5,-97</position>
<input>
<ID>IN_0</ID>838 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>466</ID>
<type>DA_FROM</type>
<position>113,-230</position>
<input>
<ID>IN_0</ID>575 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>856</ID>
<type>DA_FROM</type>
<position>370.5,-99.5</position>
<input>
<ID>IN_0</ID>839 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>857</ID>
<type>DA_FROM</type>
<position>371,-102.5</position>
<input>
<ID>IN_0</ID>840 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>468</ID>
<type>DA_FROM</type>
<position>113,-232.5</position>
<input>
<ID>IN_0</ID>576 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>858</ID>
<type>DA_FROM</type>
<position>371,-105</position>
<input>
<ID>IN_0</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>859</ID>
<type>DE_TO</type>
<position>399.5,-93.5</position>
<input>
<ID>IN_0</ID>842 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load-ADREG</lparam></gate>
<gate>
<ID>470</ID>
<type>DE_TO</type>
<position>141.5,-221</position>
<input>
<ID>IN_0</ID>577 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Res-Acc</lparam></gate>
<gate>
<ID>860</ID>
<type>DE_OR8</type>
<position>393,-159.5</position>
<input>
<ID>IN_0</ID>843 </input>
<input>
<ID>IN_1</ID>844 </input>
<input>
<ID>IN_2</ID>845 </input>
<input>
<ID>IN_3</ID>846 </input>
<input>
<ID>IN_4</ID>850 </input>
<input>
<ID>IN_5</ID>849 </input>
<input>
<ID>IN_6</ID>848 </input>
<input>
<ID>IN_7</ID>847 </input>
<output>
<ID>OUT</ID>851 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>861</ID>
<type>DA_FROM</type>
<position>383,-152.5</position>
<input>
<ID>IN_0</ID>843 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>862</ID>
<type>DA_FROM</type>
<position>375,-155</position>
<input>
<ID>IN_0</ID>844 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>863</ID>
<type>DA_FROM</type>
<position>373.5,-157.5</position>
<input>
<ID>IN_0</ID>845 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>864</ID>
<type>DA_FROM</type>
<position>373.5,-160</position>
<input>
<ID>IN_0</ID>846 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>865</ID>
<type>DA_FROM</type>
<position>373.5,-163</position>
<input>
<ID>IN_0</ID>847 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>866</ID>
<type>DA_FROM</type>
<position>373.5,-165.5</position>
<input>
<ID>IN_0</ID>848 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>867</ID>
<type>DA_FROM</type>
<position>374,-168.5</position>
<input>
<ID>IN_0</ID>849 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>868</ID>
<type>DA_FROM</type>
<position>374,-171</position>
<input>
<ID>IN_0</ID>850 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>869</ID>
<type>DE_TO</type>
<position>402.5,-159.5</position>
<input>
<ID>IN_0</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RES-ADREG</lparam></gate>
<gate>
<ID>875</ID>
<type>DE_OR8</type>
<position>393,-185.5</position>
<input>
<ID>IN_0</ID>852 </input>
<input>
<ID>IN_1</ID>853 </input>
<input>
<ID>IN_2</ID>854 </input>
<input>
<ID>IN_3</ID>855 </input>
<input>
<ID>IN_4</ID>859 </input>
<input>
<ID>IN_5</ID>858 </input>
<input>
<ID>IN_6</ID>857 </input>
<input>
<ID>IN_7</ID>856 </input>
<output>
<ID>OUT</ID>860 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>876</ID>
<type>DA_FROM</type>
<position>383,-178.5</position>
<input>
<ID>IN_0</ID>852 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>877</ID>
<type>DA_FROM</type>
<position>375,-181</position>
<input>
<ID>IN_0</ID>853 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>878</ID>
<type>DA_FROM</type>
<position>373.5,-183.5</position>
<input>
<ID>IN_0</ID>854 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>879</ID>
<type>DA_FROM</type>
<position>373.5,-186</position>
<input>
<ID>IN_0</ID>855 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>880</ID>
<type>DA_FROM</type>
<position>373.5,-189</position>
<input>
<ID>IN_0</ID>856 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>881</ID>
<type>DA_FROM</type>
<position>373.5,-191.5</position>
<input>
<ID>IN_0</ID>857 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>882</ID>
<type>DA_FROM</type>
<position>374,-194.5</position>
<input>
<ID>IN_0</ID>858 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>883</ID>
<type>DA_FROM</type>
<position>374,-197</position>
<input>
<ID>IN_0</ID>859 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>884</ID>
<type>DE_TO</type>
<position>402.5,-185.5</position>
<input>
<ID>IN_0</ID>860 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADREG-BUS</lparam></gate>
<gate>
<ID>886</ID>
<type>DE_OR8</type>
<position>390,-215.5</position>
<input>
<ID>IN_0</ID>861 </input>
<input>
<ID>IN_1</ID>862 </input>
<input>
<ID>IN_2</ID>863 </input>
<input>
<ID>IN_3</ID>864 </input>
<input>
<ID>IN_4</ID>868 </input>
<input>
<ID>IN_5</ID>867 </input>
<input>
<ID>IN_6</ID>866 </input>
<input>
<ID>IN_7</ID>865 </input>
<output>
<ID>OUT</ID>869 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>887</ID>
<type>DA_FROM</type>
<position>380,-208.5</position>
<input>
<ID>IN_0</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STA</lparam></gate>
<gate>
<ID>888</ID>
<type>DA_FROM</type>
<position>372,-211</position>
<input>
<ID>IN_0</ID>862 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STA+</lparam></gate>
<gate>
<ID>889</ID>
<type>DA_FROM</type>
<position>370.5,-213.5</position>
<input>
<ID>IN_0</ID>863 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>890</ID>
<type>DA_FROM</type>
<position>370.5,-216</position>
<input>
<ID>IN_0</ID>864 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>891</ID>
<type>DA_FROM</type>
<position>370.5,-219</position>
<input>
<ID>IN_0</ID>865 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>892</ID>
<type>DA_FROM</type>
<position>370.5,-221.5</position>
<input>
<ID>IN_0</ID>866 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>893</ID>
<type>DA_FROM</type>
<position>371,-224.5</position>
<input>
<ID>IN_0</ID>867 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>894</ID>
<type>DA_FROM</type>
<position>371,-227</position>
<input>
<ID>IN_0</ID>868 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>895</ID>
<type>DE_TO</type>
<position>399.5,-215.5</position>
<input>
<ID>IN_0</ID>869 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADREG-ADDR</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>12,-44.5</position>
<gparam>LABEL_TEXT Register Load</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>DE_OR8</type>
<position>33.5,-99.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>195 </input>
<input>
<ID>IN_2</ID>196 </input>
<input>
<ID>IN_3</ID>197 </input>
<input>
<ID>IN_4</ID>201 </input>
<input>
<ID>IN_5</ID>200 </input>
<input>
<ID>IN_6</ID>199 </input>
<input>
<ID>IN_7</ID>198 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>119</ID>
<type>DA_FROM</type>
<position>23.5,-92.5</position>
<input>
<ID>IN_0</ID>194 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADDI</lparam></gate>
<gate>
<ID>121</ID>
<type>DA_FROM</type>
<position>15.5,-95</position>
<input>
<ID>IN_0</ID>195 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MOVEI</lparam></gate>
<gate>
<ID>900</ID>
<type>DE_OR8</type>
<position>467.5,-125.5</position>
<input>
<ID>IN_0</ID>763 </input>
<input>
<ID>IN_1</ID>871 </input>
<input>
<ID>IN_2</ID>872 </input>
<input>
<ID>IN_3</ID>873 </input>
<input>
<ID>IN_4</ID>877 </input>
<input>
<ID>IN_5</ID>876 </input>
<input>
<ID>IN_6</ID>875 </input>
<input>
<ID>IN_7</ID>874 </input>
<output>
<ID>OUT</ID>878 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>14,-97.5</position>
<input>
<ID>IN_0</ID>196 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MOVE</lparam></gate>
<gate>
<ID>124</ID>
<type>DA_FROM</type>
<position>14,-100</position>
<input>
<ID>IN_0</ID>197 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>14,-103</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>127</ID>
<type>DA_FROM</type>
<position>14,-105.5</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>14.5,-108.5</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>144</ID>
<type>DA_FROM</type>
<position>14.5,-111</position>
<input>
<ID>IN_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>149</ID>
<type>DE_TO</type>
<position>43,-99.5</position>
<input>
<ID>IN_0</ID>202 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD Acc</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>52,-6</position>
<gparam>LABEL_TEXT Decode stage 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>DE_OR8</type>
<position>131,-63.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>131 </input>
<input>
<ID>IN_2</ID>133 </input>
<input>
<ID>IN_3</ID>134 </input>
<input>
<ID>IN_4</ID>138 </input>
<input>
<ID>IN_5</ID>137 </input>
<input>
<ID>IN_6</ID>136 </input>
<input>
<ID>IN_7</ID>135 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>154</ID>
<type>DA_FROM</type>
<position>121,-56.5</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MOVE</lparam></gate>
<gate>
<ID>935</ID>
<type>DE_OR8</type>
<position>389.5,-240</position>
<input>
<ID>IN_0</ID>905 </input>
<input>
<ID>IN_1</ID>906 </input>
<input>
<ID>IN_2</ID>907 </input>
<input>
<ID>IN_3</ID>908 </input>
<input>
<ID>IN_4</ID>912 </input>
<input>
<ID>IN_5</ID>911 </input>
<input>
<ID>IN_6</ID>910 </input>
<input>
<ID>IN_7</ID>909 </input>
<output>
<ID>OUT</ID>913 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>157</ID>
<type>DA_FROM</type>
<position>113,-59</position>
<input>
<ID>IN_0</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STORE</lparam></gate>
<gate>
<ID>936</ID>
<type>DA_FROM</type>
<position>379.5,-233</position>
<input>
<ID>IN_0</ID>905 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>937</ID>
<type>DA_FROM</type>
<position>371.5,-235.5</position>
<input>
<ID>IN_0</ID>906 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>159</ID>
<type>DE_TO</type>
<position>34,-3</position>
<input>
<ID>IN_0</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>938</ID>
<type>DA_FROM</type>
<position>370,-238</position>
<input>
<ID>IN_0</ID>907 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>939</ID>
<type>DA_FROM</type>
<position>370,-240.5</position>
<input>
<ID>IN_0</ID>908 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>161</ID>
<type>FF_GND</type>
<position>30.5,-3</position>
<output>
<ID>OUT_0</ID>132 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>940</ID>
<type>DA_FROM</type>
<position>370,-243.5</position>
<input>
<ID>IN_0</ID>909 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>162</ID>
<type>DA_FROM</type>
<position>111.5,-61.5</position>
<input>
<ID>IN_0</ID>133 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>941</ID>
<type>DA_FROM</type>
<position>370,-246</position>
<input>
<ID>IN_0</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>163</ID>
<type>DA_FROM</type>
<position>111.5,-64</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>942</ID>
<type>DA_FROM</type>
<position>370.5,-249</position>
<input>
<ID>IN_0</ID>911 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>164</ID>
<type>DA_FROM</type>
<position>111.5,-67</position>
<input>
<ID>IN_0</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>943</ID>
<type>DA_FROM</type>
<position>370.5,-251.5</position>
<input>
<ID>IN_0</ID>912 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>111.5,-69.5</position>
<input>
<ID>IN_0</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>944</ID>
<type>DE_TO</type>
<position>399,-240</position>
<input>
<ID>IN_0</ID>913 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Res-ADDR</lparam></gate>
<gate>
<ID>166</ID>
<type>DA_FROM</type>
<position>112,-72.5</position>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>167</ID>
<type>DA_FROM</type>
<position>112,-75</position>
<input>
<ID>IN_0</ID>138 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>168</ID>
<type>DE_OR8</type>
<position>325,-65</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>204 </input>
<input>
<ID>IN_2</ID>205 </input>
<input>
<ID>IN_3</ID>206 </input>
<input>
<ID>IN_4</ID>210 </input>
<input>
<ID>IN_5</ID>209 </input>
<input>
<ID>IN_6</ID>208 </input>
<input>
<ID>IN_7</ID>207 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>947</ID>
<type>DA_FROM</type>
<position>457.5,-118.5</position>
<input>
<ID>IN_0</ID>763 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>169</ID>
<type>DE_TO</type>
<position>140.5,-63.5</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-AD</lparam></gate>
<gate>
<ID>170</ID>
<type>DE_OR8</type>
<position>132,-91.5</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>141 </input>
<input>
<ID>IN_2</ID>142 </input>
<input>
<ID>IN_3</ID>143 </input>
<input>
<ID>IN_4</ID>147 </input>
<input>
<ID>IN_5</ID>146 </input>
<input>
<ID>IN_6</ID>145 </input>
<input>
<ID>IN_7</ID>144 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>171</ID>
<type>DA_FROM</type>
<position>122,-84.5</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADDI</lparam></gate>
<gate>
<ID>172</ID>
<type>DA_FROM</type>
<position>114,-87</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MOVEI</lparam></gate>
<gate>
<ID>173</ID>
<type>DA_FROM</type>
<position>112.5,-89.5</position>
<input>
<ID>IN_0</ID>142 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>174</ID>
<type>DA_FROM</type>
<position>112.5,-92</position>
<input>
<ID>IN_0</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>175</ID>
<type>DA_FROM</type>
<position>112.5,-95</position>
<input>
<ID>IN_0</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>176</ID>
<type>DA_FROM</type>
<position>112.5,-97.5</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>177</ID>
<type>DA_FROM</type>
<position>113,-100.5</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>113,-103</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>179</ID>
<type>DE_TO</type>
<position>141.5,-91.5</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Imm</lparam></gate>
<gate>
<ID>180</ID>
<type>DE_OR8</type>
<position>33.5,-136</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>150 </input>
<input>
<ID>IN_2</ID>151 </input>
<input>
<ID>IN_3</ID>152 </input>
<input>
<ID>IN_4</ID>156 </input>
<input>
<ID>IN_5</ID>155 </input>
<input>
<ID>IN_6</ID>154 </input>
<input>
<ID>IN_7</ID>153 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>181</ID>
<type>DA_FROM</type>
<position>23.5,-129</position>
<input>
<ID>IN_0</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STORE</lparam></gate>
<gate>
<ID>182</ID>
<type>DA_FROM</type>
<position>15.5,-131.5</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STA</lparam></gate>
<gate>
<ID>961</ID>
<type>DA_FROM</type>
<position>449.5,-121</position>
<input>
<ID>IN_0</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>183</ID>
<type>DA_FROM</type>
<position>14,-134</position>
<input>
<ID>IN_0</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STA+</lparam></gate>
<gate>
<ID>184</ID>
<type>DA_FROM</type>
<position>14,-136.5</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>185</ID>
<type>DA_FROM</type>
<position>14,-139.5</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>186</ID>
<type>DA_FROM</type>
<position>14,-142</position>
<input>
<ID>IN_0</ID>154 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>187</ID>
<type>DA_FROM</type>
<position>14.5,-145</position>
<input>
<ID>IN_0</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>188</ID>
<type>DA_FROM</type>
<position>14.5,-147.5</position>
<input>
<ID>IN_0</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>189</ID>
<type>DE_TO</type>
<position>43,-136</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Mem Write</lparam></gate>
<gate>
<ID>190</ID>
<type>DE_OR8</type>
<position>134,-129.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>159 </input>
<input>
<ID>IN_2</ID>160 </input>
<input>
<ID>IN_3</ID>161 </input>
<input>
<ID>IN_4</ID>165 </input>
<input>
<ID>IN_5</ID>164 </input>
<input>
<ID>IN_6</ID>163 </input>
<input>
<ID>IN_7</ID>162 </input>
<output>
<ID>OUT</ID>166 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>579</ID>
<type>DE_OR8</type>
<position>173,-90</position>
<input>
<ID>IN_0</ID>705 </input>
<input>
<ID>IN_1</ID>706 </input>
<input>
<ID>IN_2</ID>707 </input>
<input>
<ID>IN_3</ID>708 </input>
<input>
<ID>IN_4</ID>712 </input>
<input>
<ID>IN_5</ID>711 </input>
<input>
<ID>IN_6</ID>710 </input>
<input>
<ID>IN_7</ID>709 </input>
<output>
<ID>OUT</ID>713 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>191</ID>
<type>DA_FROM</type>
<position>124,-122.5</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>969</ID>
<type>DA_FROM</type>
<position>448,-123.5</position>
<input>
<ID>IN_0</ID>872 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>580</ID>
<type>DA_FROM</type>
<position>163,-83</position>
<input>
<ID>IN_0</ID>705 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADDI</lparam></gate>
<gate>
<ID>192</ID>
<type>DA_FROM</type>
<position>116,-125</position>
<input>
<ID>IN_0</ID>159 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MOVE</lparam></gate>
<gate>
<ID>581</ID>
<type>DA_FROM</type>
<position>155,-85.5</position>
<input>
<ID>IN_0</ID>706 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>582</ID>
<type>DA_FROM</type>
<position>153.5,-88</position>
<input>
<ID>IN_0</ID>707 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>193</ID>
<type>DA_FROM</type>
<position>114.5,-127.5</position>
<input>
<ID>IN_0</ID>160 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>583</ID>
<type>DA_FROM</type>
<position>153.5,-90.5</position>
<input>
<ID>IN_0</ID>708 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>194</ID>
<type>DA_FROM</type>
<position>114.5,-130</position>
<input>
<ID>IN_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>584</ID>
<type>DA_FROM</type>
<position>153.5,-93.5</position>
<input>
<ID>IN_0</ID>709 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>195</ID>
<type>DA_FROM</type>
<position>114.5,-133</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>585</ID>
<type>DA_FROM</type>
<position>153.5,-96</position>
<input>
<ID>IN_0</ID>710 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>196</ID>
<type>DA_FROM</type>
<position>114.5,-135.5</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>197</ID>
<type>DA_FROM</type>
<position>115,-138.5</position>
<input>
<ID>IN_0</ID>164 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>587</ID>
<type>DA_FROM</type>
<position>154,-99</position>
<input>
<ID>IN_0</ID>711 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>198</ID>
<type>DA_FROM</type>
<position>115,-141</position>
<input>
<ID>IN_0</ID>165 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>199</ID>
<type>DE_TO</type>
<position>143.5,-129.5</position>
<input>
<ID>IN_0</ID>166 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Mem Read</lparam></gate>
<gate>
<ID>200</ID>
<type>DA_FROM</type>
<position>315,-58</position>
<input>
<ID>IN_0</ID>203 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BRA</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_LABEL</type>
<position>107.5,-44.5</position>
<gparam>LABEL_TEXT Bus and Memory Controls</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>DA_FROM</type>
<position>307,-60.5</position>
<input>
<ID>IN_0</ID>204 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>981</ID>
<type>DA_FROM</type>
<position>448,-126</position>
<input>
<ID>IN_0</ID>873 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>982</ID>
<type>DA_FROM</type>
<position>448,-129</position>
<input>
<ID>IN_0</ID>874 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>204</ID>
<type>DA_FROM</type>
<position>305.5,-63</position>
<input>
<ID>IN_0</ID>205 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>983</ID>
<type>DA_FROM</type>
<position>448,-131.5</position>
<input>
<ID>IN_0</ID>875 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>205</ID>
<type>DA_FROM</type>
<position>305.5,-65.5</position>
<input>
<ID>IN_0</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>595</ID>
<type>DA_FROM</type>
<position>154,-101.5</position>
<input>
<ID>IN_0</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>206</ID>
<type>DA_FROM</type>
<position>305.5,-68.5</position>
<input>
<ID>IN_0</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>985</ID>
<type>DA_FROM</type>
<position>448.5,-134.5</position>
<input>
<ID>IN_0</ID>876 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>207</ID>
<type>DA_FROM</type>
<position>305.5,-71</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>208</ID>
<type>DA_FROM</type>
<position>306,-74</position>
<input>
<ID>IN_0</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>987</ID>
<type>DA_FROM</type>
<position>448.5,-137</position>
<input>
<ID>IN_0</ID>877 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>598</ID>
<type>DE_TO</type>
<position>182.5,-90</position>
<input>
<ID>IN_0</ID>713 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID StatEn</lparam></gate>
<gate>
<ID>209</ID>
<type>DA_FROM</type>
<position>306,-76.5</position>
<input>
<ID>IN_0</ID>210 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>210</ID>
<type>DE_TO</type>
<position>334.5,-65</position>
<input>
<ID>IN_0</ID>211 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC EXS</lparam></gate>
<gate>
<ID>989</ID>
<type>DE_TO</type>
<position>477,-125.5</position>
<input>
<ID>IN_0</ID>878 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BUS-SP</lparam></gate>
<gate>
<ID>211</ID>
<type>DE_OR8</type>
<position>33.5,-66.5</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>168 </input>
<input>
<ID>IN_2</ID>169 </input>
<input>
<ID>IN_3</ID>170 </input>
<input>
<ID>IN_4</ID>174 </input>
<input>
<ID>IN_5</ID>173 </input>
<input>
<ID>IN_6</ID>172 </input>
<input>
<ID>IN_7</ID>171 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>212</ID>
<type>DA_FROM</type>
<position>23.5,-59.5</position>
<input>
<ID>IN_0</ID>167 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID JMP</lparam></gate>
<gate>
<ID>991</ID>
<type>DE_OR8</type>
<position>465,-59.5</position>
<input>
<ID>IN_0</ID>902 </input>
<input>
<ID>IN_1</ID>914 </input>
<input>
<ID>IN_2</ID>915 </input>
<input>
<ID>IN_3</ID>916 </input>
<input>
<ID>IN_4</ID>1006 </input>
<input>
<ID>IN_5</ID>1005 </input>
<input>
<ID>IN_6</ID>1004 </input>
<input>
<ID>IN_7</ID>917 </input>
<output>
<ID>OUT</ID>1007 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>213</ID>
<type>DA_FROM</type>
<position>15.5,-62</position>
<input>
<ID>IN_0</ID>168 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BRA</lparam></gate>
<gate>
<ID>214</ID>
<type>DA_FROM</type>
<position>14,-64.5</position>
<input>
<ID>IN_0</ID>169 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>993</ID>
<type>DA_FROM</type>
<position>455,-52.5</position>
<input>
<ID>IN_0</ID>902 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>215</ID>
<type>DA_FROM</type>
<position>14,-67</position>
<input>
<ID>IN_0</ID>170 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>216</ID>
<type>DA_FROM</type>
<position>14,-70</position>
<input>
<ID>IN_0</ID>171 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>995</ID>
<type>DA_FROM</type>
<position>447,-55</position>
<input>
<ID>IN_0</ID>914 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>217</ID>
<type>DA_FROM</type>
<position>14,-72.5</position>
<input>
<ID>IN_0</ID>172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>218</ID>
<type>DA_FROM</type>
<position>14.5,-75.5</position>
<input>
<ID>IN_0</ID>173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>997</ID>
<type>DA_FROM</type>
<position>445.5,-57.5</position>
<input>
<ID>IN_0</ID>915 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>219</ID>
<type>DA_FROM</type>
<position>14.5,-78</position>
<input>
<ID>IN_0</ID>174 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>220</ID>
<type>DE_TO</type>
<position>43,-66.5</position>
<input>
<ID>IN_0</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load PC</lparam></gate>
<gate>
<ID>610</ID>
<type>DE_OR8</type>
<position>233.5,-129.5</position>
<input>
<ID>IN_0</ID>538 </input>
<input>
<ID>IN_1</ID>539 </input>
<input>
<ID>IN_2</ID>540 </input>
<input>
<ID>IN_3</ID>541 </input>
<input>
<ID>IN_4</ID>545 </input>
<input>
<ID>IN_5</ID>544 </input>
<input>
<ID>IN_6</ID>543 </input>
<input>
<ID>IN_7</ID>542 </input>
<output>
<ID>OUT</ID>546 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>221</ID>
<type>DE_OR8</type>
<position>324.5,-91.5</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>213 </input>
<input>
<ID>IN_2</ID>214 </input>
<input>
<ID>IN_3</ID>215 </input>
<input>
<ID>IN_4</ID>219 </input>
<input>
<ID>IN_5</ID>218 </input>
<input>
<ID>IN_6</ID>217 </input>
<input>
<ID>IN_7</ID>216 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1000</ID>
<type>DA_FROM</type>
<position>445.5,-60</position>
<input>
<ID>IN_0</ID>916 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>611</ID>
<type>DA_FROM</type>
<position>223.5,-122.5</position>
<input>
<ID>IN_0</ID>538 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>222</ID>
<type>DA_FROM</type>
<position>314.5,-84.5</position>
<input>
<ID>IN_0</ID>212 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BRA</lparam></gate>
<gate>
<ID>612</ID>
<type>DA_FROM</type>
<position>215.5,-125</position>
<input>
<ID>IN_0</ID>539 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>223</ID>
<type>DA_FROM</type>
<position>306.5,-87</position>
<input>
<ID>IN_0</ID>213 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID JMP</lparam></gate>
<gate>
<ID>1002</ID>
<type>DA_FROM</type>
<position>445.5,-63</position>
<input>
<ID>IN_0</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>613</ID>
<type>DA_FROM</type>
<position>214,-127.5</position>
<input>
<ID>IN_0</ID>540 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>224</ID>
<type>DA_FROM</type>
<position>305,-89.5</position>
<input>
<ID>IN_0</ID>214 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1003</ID>
<type>DA_FROM</type>
<position>445.5,-65.5</position>
<input>
<ID>IN_0</ID>1004 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>614</ID>
<type>DA_FROM</type>
<position>214,-130</position>
<input>
<ID>IN_0</ID>541 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>225</ID>
<type>DA_FROM</type>
<position>305,-92</position>
<input>
<ID>IN_0</ID>215 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1004</ID>
<type>DA_FROM</type>
<position>446,-68.5</position>
<input>
<ID>IN_0</ID>1005 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>615</ID>
<type>DA_FROM</type>
<position>214,-133</position>
<input>
<ID>IN_0</ID>542 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>226</ID>
<type>DA_FROM</type>
<position>305,-95</position>
<input>
<ID>IN_0</ID>216 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1005</ID>
<type>DA_FROM</type>
<position>446,-71</position>
<input>
<ID>IN_0</ID>1006 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>616</ID>
<type>DA_FROM</type>
<position>214,-135.5</position>
<input>
<ID>IN_0</ID>543 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>227</ID>
<type>DA_FROM</type>
<position>305,-97.5</position>
<input>
<ID>IN_0</ID>217 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1006</ID>
<type>DE_TO</type>
<position>474.5,-59.5</position>
<input>
<ID>IN_0</ID>1007 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INC-SP</lparam></gate>
<gate>
<ID>617</ID>
<type>DA_FROM</type>
<position>214.5,-138.5</position>
<input>
<ID>IN_0</ID>544 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>228</ID>
<type>DA_FROM</type>
<position>305.5,-100.5</position>
<input>
<ID>IN_0</ID>218 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1007</ID>
<type>DE_OR8</type>
<position>465,-91</position>
<input>
<ID>IN_0</ID>1008 </input>
<input>
<ID>IN_1</ID>1009 </input>
<input>
<ID>IN_2</ID>1010 </input>
<input>
<ID>IN_3</ID>1011 </input>
<input>
<ID>IN_4</ID>1015 </input>
<input>
<ID>IN_5</ID>1014 </input>
<input>
<ID>IN_6</ID>1013 </input>
<input>
<ID>IN_7</ID>1012 </input>
<output>
<ID>OUT</ID>1016 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>618</ID>
<type>DA_FROM</type>
<position>214.5,-141</position>
<input>
<ID>IN_0</ID>545 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>229</ID>
<type>DA_FROM</type>
<position>305.5,-103</position>
<input>
<ID>IN_0</ID>219 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1008</ID>
<type>DA_FROM</type>
<position>455,-84</position>
<input>
<ID>IN_0</ID>1008 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>619</ID>
<type>DE_TO</type>
<position>243,-129.5</position>
<input>
<ID>IN_0</ID>546 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZero</lparam></gate>
<gate>
<ID>230</ID>
<type>DE_TO</type>
<position>334,-91.5</position>
<input>
<ID>IN_0</ID>220 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-PC</lparam></gate>
<gate>
<ID>1009</ID>
<type>DA_FROM</type>
<position>447,-86.5</position>
<input>
<ID>IN_0</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>231</ID>
<type>DE_OR8</type>
<position>326,-123.5</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>222 </input>
<input>
<ID>IN_2</ID>223 </input>
<input>
<ID>IN_3</ID>224 </input>
<input>
<ID>IN_4</ID>228 </input>
<input>
<ID>IN_5</ID>227 </input>
<input>
<ID>IN_6</ID>226 </input>
<input>
<ID>IN_7</ID>225 </input>
<output>
<ID>OUT</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1010</ID>
<type>DA_FROM</type>
<position>445.5,-89</position>
<input>
<ID>IN_0</ID>1010 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>621</ID>
<type>AA_LABEL</type>
<position>220,-43</position>
<gparam>LABEL_TEXT ALU Controls</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>DA_FROM</type>
<position>312.5,-116</position>
<input>
<ID>IN_0</ID>221 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1011</ID>
<type>DA_FROM</type>
<position>445.5,-91.5</position>
<input>
<ID>IN_0</ID>1011 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>622</ID>
<type>DE_OR8</type>
<position>231,-63.5</position>
<input>
<ID>IN_0</ID>547 </input>
<input>
<ID>IN_1</ID>548 </input>
<input>
<ID>IN_2</ID>549 </input>
<input>
<ID>IN_3</ID>550 </input>
<input>
<ID>IN_4</ID>554 </input>
<input>
<ID>IN_5</ID>553 </input>
<input>
<ID>IN_6</ID>552 </input>
<input>
<ID>IN_7</ID>551 </input>
<output>
<ID>OUT</ID>555 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>233</ID>
<type>DA_FROM</type>
<position>308,-119</position>
<input>
<ID>IN_0</ID>222 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID JMP</lparam></gate>
<gate>
<ID>1012</ID>
<type>DA_FROM</type>
<position>445.5,-94.5</position>
<input>
<ID>IN_0</ID>1012 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>623</ID>
<type>DA_FROM</type>
<position>221,-56.5</position>
<input>
<ID>IN_0</ID>547 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>234</ID>
<type>DA_FROM</type>
<position>306.5,-121.5</position>
<input>
<ID>IN_0</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1013</ID>
<type>DA_FROM</type>
<position>445.5,-97</position>
<input>
<ID>IN_0</ID>1013 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>624</ID>
<type>DA_FROM</type>
<position>213,-59</position>
<input>
<ID>IN_0</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>235</ID>
<type>DA_FROM</type>
<position>306.5,-124</position>
<input>
<ID>IN_0</ID>224 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1014</ID>
<type>DA_FROM</type>
<position>446,-100</position>
<input>
<ID>IN_0</ID>1014 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>625</ID>
<type>DA_FROM</type>
<position>211.5,-61.5</position>
<input>
<ID>IN_0</ID>549 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>236</ID>
<type>DA_FROM</type>
<position>306.5,-127</position>
<input>
<ID>IN_0</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1015</ID>
<type>DA_FROM</type>
<position>446,-102.5</position>
<input>
<ID>IN_0</ID>1015 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>626</ID>
<type>DA_FROM</type>
<position>211.5,-64</position>
<input>
<ID>IN_0</ID>550 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>237</ID>
<type>DA_FROM</type>
<position>306.5,-129.5</position>
<input>
<ID>IN_0</ID>226 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1016</ID>
<type>DE_TO</type>
<position>474.5,-91</position>
<input>
<ID>IN_0</ID>1016 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load-SP</lparam></gate>
<gate>
<ID>627</ID>
<type>DA_FROM</type>
<position>211.5,-67</position>
<input>
<ID>IN_0</ID>551 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>238</ID>
<type>DA_FROM</type>
<position>307,-132.5</position>
<input>
<ID>IN_0</ID>227 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1017</ID>
<type>DE_OR8</type>
<position>468,-157</position>
<input>
<ID>IN_0</ID>1017 </input>
<input>
<ID>IN_1</ID>1018 </input>
<input>
<ID>IN_2</ID>1019 </input>
<input>
<ID>IN_3</ID>1020 </input>
<input>
<ID>IN_4</ID>1024 </input>
<input>
<ID>IN_5</ID>1023 </input>
<input>
<ID>IN_6</ID>1022 </input>
<input>
<ID>IN_7</ID>1021 </input>
<output>
<ID>OUT</ID>1025 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>628</ID>
<type>DA_FROM</type>
<position>211.5,-69.5</position>
<input>
<ID>IN_0</ID>552 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>239</ID>
<type>DA_FROM</type>
<position>307,-135</position>
<input>
<ID>IN_0</ID>228 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1018</ID>
<type>DA_FROM</type>
<position>458,-150</position>
<input>
<ID>IN_0</ID>1017 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>629</ID>
<type>DA_FROM</type>
<position>212,-72.5</position>
<input>
<ID>IN_0</ID>553 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>240</ID>
<type>DE_TO</type>
<position>335.5,-123.5</position>
<input>
<ID>IN_0</ID>229 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCDIR</lparam></gate>
<gate>
<ID>1019</ID>
<type>DA_FROM</type>
<position>450,-152.5</position>
<input>
<ID>IN_0</ID>1018 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>630</ID>
<type>DA_FROM</type>
<position>212,-75</position>
<input>
<ID>IN_0</ID>554 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>241</ID>
<type>AA_LABEL</type>
<position>301,-40.5</position>
<gparam>LABEL_TEXT PC Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1020</ID>
<type>DA_FROM</type>
<position>448.5,-155</position>
<input>
<ID>IN_0</ID>1019 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>631</ID>
<type>DE_TO</type>
<position>240.5,-63.5</position>
<input>
<ID>IN_0</ID>555 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUBA</lparam></gate>
<gate>
<ID>242</ID>
<type>DE_OR8</type>
<position>325.5,-146</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>231 </input>
<input>
<ID>IN_2</ID>232 </input>
<input>
<ID>IN_3</ID>233 </input>
<input>
<ID>IN_4</ID>237 </input>
<input>
<ID>IN_5</ID>236 </input>
<input>
<ID>IN_6</ID>235 </input>
<input>
<ID>IN_7</ID>234 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1021</ID>
<type>DA_FROM</type>
<position>448.5,-157.5</position>
<input>
<ID>IN_0</ID>1020 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>243</ID>
<type>DA_FROM</type>
<position>315.5,-139</position>
<input>
<ID>IN_0</ID>230 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BRA</lparam></gate>
<gate>
<ID>1022</ID>
<type>DA_FROM</type>
<position>448.5,-160.5</position>
<input>
<ID>IN_0</ID>1021 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>633</ID>
<type>DE_OR8</type>
<position>231,-95</position>
<input>
<ID>IN_0</ID>556 </input>
<input>
<ID>IN_1</ID>557 </input>
<input>
<ID>IN_2</ID>558 </input>
<input>
<ID>IN_3</ID>559 </input>
<input>
<ID>IN_4</ID>563 </input>
<input>
<ID>IN_5</ID>562 </input>
<input>
<ID>IN_6</ID>561 </input>
<input>
<ID>IN_7</ID>560 </input>
<output>
<ID>OUT</ID>564 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>244</ID>
<type>DA_FROM</type>
<position>307.5,-141.5</position>
<input>
<ID>IN_0</ID>231 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1023</ID>
<type>DA_FROM</type>
<position>448.5,-163</position>
<input>
<ID>IN_0</ID>1022 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>634</ID>
<type>DA_FROM</type>
<position>221,-88</position>
<input>
<ID>IN_0</ID>556 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>245</ID>
<type>DA_FROM</type>
<position>306,-144</position>
<input>
<ID>IN_0</ID>232 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1024</ID>
<type>DA_FROM</type>
<position>449,-166</position>
<input>
<ID>IN_0</ID>1023 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>635</ID>
<type>DA_FROM</type>
<position>213,-90.5</position>
<input>
<ID>IN_0</ID>557 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>246</ID>
<type>DA_FROM</type>
<position>306,-146.5</position>
<input>
<ID>IN_0</ID>233 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1025</ID>
<type>DA_FROM</type>
<position>449,-168.5</position>
<input>
<ID>IN_0</ID>1024 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>636</ID>
<type>DA_FROM</type>
<position>211.5,-93</position>
<input>
<ID>IN_0</ID>558 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>247</ID>
<type>DA_FROM</type>
<position>306,-149.5</position>
<input>
<ID>IN_0</ID>234 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1026</ID>
<type>DE_TO</type>
<position>477.5,-157</position>
<input>
<ID>IN_0</ID>1025 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RES-SP</lparam></gate>
<gate>
<ID>637</ID>
<type>DA_FROM</type>
<position>211.5,-95.5</position>
<input>
<ID>IN_0</ID>559 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>248</ID>
<type>DA_FROM</type>
<position>306,-152</position>
<input>
<ID>IN_0</ID>235 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1027</ID>
<type>DE_OR8</type>
<position>468,-183</position>
<input>
<ID>IN_0</ID>1026 </input>
<input>
<ID>IN_1</ID>1027 </input>
<input>
<ID>IN_2</ID>1028 </input>
<input>
<ID>IN_3</ID>1029 </input>
<input>
<ID>IN_4</ID>1033 </input>
<input>
<ID>IN_5</ID>1032 </input>
<input>
<ID>IN_6</ID>1031 </input>
<input>
<ID>IN_7</ID>1030 </input>
<output>
<ID>OUT</ID>1034 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>638</ID>
<type>DA_FROM</type>
<position>211.5,-98.5</position>
<input>
<ID>IN_0</ID>560 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>249</ID>
<type>DA_FROM</type>
<position>306.5,-155</position>
<input>
<ID>IN_0</ID>236 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1028</ID>
<type>DA_FROM</type>
<position>458,-176</position>
<input>
<ID>IN_0</ID>1026 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>639</ID>
<type>DA_FROM</type>
<position>211.5,-101</position>
<input>
<ID>IN_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>250</ID>
<type>DA_FROM</type>
<position>306.5,-157.5</position>
<input>
<ID>IN_0</ID>237 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1029</ID>
<type>DA_FROM</type>
<position>450,-178.5</position>
<input>
<ID>IN_0</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>640</ID>
<type>DA_FROM</type>
<position>212,-104</position>
<input>
<ID>IN_0</ID>562 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>251</ID>
<type>DE_TO</type>
<position>335,-146</position>
<input>
<ID>IN_0</ID>238 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Offset</lparam></gate>
<gate>
<ID>1030</ID>
<type>DA_FROM</type>
<position>448.5,-181</position>
<input>
<ID>IN_0</ID>1028 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>641</ID>
<type>DA_FROM</type>
<position>212,-106.5</position>
<input>
<ID>IN_0</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>252</ID>
<type>DE_OR8</type>
<position>131,-191</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>240 </input>
<input>
<ID>IN_2</ID>241 </input>
<input>
<ID>IN_3</ID>242 </input>
<input>
<ID>IN_4</ID>246 </input>
<input>
<ID>IN_5</ID>245 </input>
<input>
<ID>IN_6</ID>244 </input>
<input>
<ID>IN_7</ID>243 </input>
<output>
<ID>OUT</ID>247 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1031</ID>
<type>DA_FROM</type>
<position>448.5,-183.5</position>
<input>
<ID>IN_0</ID>1029 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>642</ID>
<type>DE_TO</type>
<position>240.5,-95</position>
<input>
<ID>IN_0</ID>564 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUBB</lparam></gate>
<gate>
<ID>253</ID>
<type>DA_FROM</type>
<position>121,-184</position>
<input>
<ID>IN_0</ID>239 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1032</ID>
<type>DA_FROM</type>
<position>448.5,-186.5</position>
<input>
<ID>IN_0</ID>1030 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>643</ID>
<type>DE_OR8</type>
<position>131,-156.5</position>
<input>
<ID>IN_0</ID>565 </input>
<input>
<ID>IN_1</ID>566 </input>
<input>
<ID>IN_2</ID>567 </input>
<input>
<ID>IN_3</ID>568 </input>
<input>
<ID>IN_4</ID>572 </input>
<input>
<ID>IN_5</ID>571 </input>
<input>
<ID>IN_6</ID>570 </input>
<input>
<ID>IN_7</ID>569 </input>
<output>
<ID>OUT</ID>573 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>254</ID>
<type>DA_FROM</type>
<position>113,-186.5</position>
<input>
<ID>IN_0</ID>240 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1033</ID>
<type>DA_FROM</type>
<position>448.5,-189</position>
<input>
<ID>IN_0</ID>1031 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>644</ID>
<type>DA_FROM</type>
<position>121,-149.5</position>
<input>
<ID>IN_0</ID>565 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STORE</lparam></gate>
<gate>
<ID>1034</ID>
<type>DA_FROM</type>
<position>449,-192</position>
<input>
<ID>IN_0</ID>1032 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>645</ID>
<type>DA_FROM</type>
<position>113,-152</position>
<input>
<ID>IN_0</ID>566 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STA</lparam></gate>
<gate>
<ID>256</ID>
<type>DA_FROM</type>
<position>111.5,-189</position>
<input>
<ID>IN_0</ID>241 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1035</ID>
<type>DA_FROM</type>
<position>449,-194.5</position>
<input>
<ID>IN_0</ID>1033 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>646</ID>
<type>DA_FROM</type>
<position>111.5,-154.5</position>
<input>
<ID>IN_0</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STA+</lparam></gate>
<gate>
<ID>257</ID>
<type>DA_FROM</type>
<position>111.5,-191.5</position>
<input>
<ID>IN_0</ID>242 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1036</ID>
<type>DE_TO</type>
<position>477.5,-183</position>
<input>
<ID>IN_0</ID>1034 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SP-BUS</lparam></gate>
<gate>
<ID>647</ID>
<type>DA_FROM</type>
<position>111.5,-157</position>
<input>
<ID>IN_0</ID>568 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>258</ID>
<type>DA_FROM</type>
<position>111.5,-194.5</position>
<input>
<ID>IN_0</ID>243 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1037</ID>
<type>DE_OR8</type>
<position>465,-213</position>
<input>
<ID>IN_0</ID>1035 </input>
<input>
<ID>IN_1</ID>1036 </input>
<input>
<ID>IN_2</ID>1037 </input>
<input>
<ID>IN_3</ID>1038 </input>
<input>
<ID>IN_4</ID>1042 </input>
<input>
<ID>IN_5</ID>1041 </input>
<input>
<ID>IN_6</ID>1040 </input>
<input>
<ID>IN_7</ID>1039 </input>
<output>
<ID>OUT</ID>1043 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>648</ID>
<type>DA_FROM</type>
<position>111.5,-160</position>
<input>
<ID>IN_0</ID>569 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>259</ID>
<type>DA_FROM</type>
<position>111.5,-197</position>
<input>
<ID>IN_0</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1038</ID>
<type>DA_FROM</type>
<position>455,-206</position>
<input>
<ID>IN_0</ID>1035 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>649</ID>
<type>DA_FROM</type>
<position>111.5,-162.5</position>
<input>
<ID>IN_0</ID>570 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>260</ID>
<type>DA_FROM</type>
<position>112,-200</position>
<input>
<ID>IN_0</ID>245 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1039</ID>
<type>DA_FROM</type>
<position>447,-208.5</position>
<input>
<ID>IN_0</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>650</ID>
<type>DA_FROM</type>
<position>112,-165.5</position>
<input>
<ID>IN_0</ID>571 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>261</ID>
<type>DA_FROM</type>
<position>112,-202.5</position>
<input>
<ID>IN_0</ID>246 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1040</ID>
<type>DA_FROM</type>
<position>445.5,-211</position>
<input>
<ID>IN_0</ID>1037 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>651</ID>
<type>DA_FROM</type>
<position>112,-168</position>
<input>
<ID>IN_0</ID>572 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>262</ID>
<type>DE_TO</type>
<position>140.5,-191</position>
<input>
<ID>IN_0</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-BUS</lparam></gate>
<gate>
<ID>1041</ID>
<type>DA_FROM</type>
<position>445.5,-213.5</position>
<input>
<ID>IN_0</ID>1038 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>652</ID>
<type>DE_TO</type>
<position>140.5,-156.5</position>
<input>
<ID>IN_0</ID>573 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Acc-Bus</lparam></gate>
<gate>
<ID>1042</ID>
<type>DA_FROM</type>
<position>445.5,-216.5</position>
<input>
<ID>IN_0</ID>1039 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1043</ID>
<type>DA_FROM</type>
<position>445.5,-219</position>
<input>
<ID>IN_0</ID>1040 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1044</ID>
<type>DA_FROM</type>
<position>446,-222</position>
<input>
<ID>IN_0</ID>1041 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1045</ID>
<type>DA_FROM</type>
<position>446,-224.5</position>
<input>
<ID>IN_0</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1046</ID>
<type>DE_TO</type>
<position>474.5,-213</position>
<input>
<ID>IN_0</ID>1043 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SP-ADDR</lparam></gate>
<gate>
<ID>1047</ID>
<type>DE_OR8</type>
<position>464.5,-237.5</position>
<input>
<ID>IN_0</ID>1044 </input>
<input>
<ID>IN_1</ID>1045 </input>
<input>
<ID>IN_2</ID>1046 </input>
<input>
<ID>IN_3</ID>1047 </input>
<input>
<ID>IN_4</ID>1051 </input>
<input>
<ID>IN_5</ID>1050 </input>
<input>
<ID>IN_6</ID>1049 </input>
<input>
<ID>IN_7</ID>1048 </input>
<output>
<ID>OUT</ID>1052 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1048</ID>
<type>DA_FROM</type>
<position>454.5,-230.5</position>
<input>
<ID>IN_0</ID>1044 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1049</ID>
<type>DA_FROM</type>
<position>446.5,-233</position>
<input>
<ID>IN_0</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1050</ID>
<type>DA_FROM</type>
<position>445,-235.5</position>
<input>
<ID>IN_0</ID>1046 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1051</ID>
<type>DA_FROM</type>
<position>445,-238</position>
<input>
<ID>IN_0</ID>1047 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1052</ID>
<type>DA_FROM</type>
<position>445,-241</position>
<input>
<ID>IN_0</ID>1048 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1053</ID>
<type>DA_FROM</type>
<position>445,-243.5</position>
<input>
<ID>IN_0</ID>1049 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1054</ID>
<type>DA_FROM</type>
<position>445.5,-246.5</position>
<input>
<ID>IN_0</ID>1050 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1055</ID>
<type>DA_FROM</type>
<position>445.5,-249</position>
<input>
<ID>IN_0</ID>1051 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1056</ID>
<type>DE_TO</type>
<position>474,-237.5</position>
<input>
<ID>IN_0</ID>1052 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Res-ADDR</lparam></gate>
<gate>
<ID>1058</ID>
<type>AA_LABEL</type>
<position>443,-39.5</position>
<gparam>LABEL_TEXT Stack</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>280</ID>
<type>DE_OR8</type>
<position>326,-168</position>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>253 </input>
<input>
<ID>IN_2</ID>254 </input>
<input>
<ID>IN_3</ID>255 </input>
<input>
<ID>IN_4</ID>259 </input>
<input>
<ID>IN_5</ID>258 </input>
<input>
<ID>IN_6</ID>257 </input>
<input>
<ID>IN_7</ID>256 </input>
<output>
<ID>OUT</ID>260 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1059</ID>
<type>DE_OR8</type>
<position>517,-59.5</position>
<input>
<ID>IN_0</ID>1053 </input>
<input>
<ID>IN_1</ID>1054 </input>
<input>
<ID>IN_2</ID>1055 </input>
<input>
<ID>IN_3</ID>1056 </input>
<input>
<ID>IN_4</ID>1060 </input>
<input>
<ID>IN_5</ID>1059 </input>
<input>
<ID>IN_6</ID>1058 </input>
<input>
<ID>IN_7</ID>1057 </input>
<output>
<ID>OUT</ID>1061 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>281</ID>
<type>DA_FROM</type>
<position>316,-161</position>
<input>
<ID>IN_0</ID>252 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1060</ID>
<type>DA_FROM</type>
<position>507,-52.5</position>
<input>
<ID>IN_0</ID>1053 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>282</ID>
<type>DA_FROM</type>
<position>308,-163.5</position>
<input>
<ID>IN_0</ID>253 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1061</ID>
<type>DA_FROM</type>
<position>499,-55</position>
<input>
<ID>IN_0</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>283</ID>
<type>DA_FROM</type>
<position>306.5,-166</position>
<input>
<ID>IN_0</ID>254 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1062</ID>
<type>DA_FROM</type>
<position>497.5,-57.5</position>
<input>
<ID>IN_0</ID>1055 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>284</ID>
<type>DA_FROM</type>
<position>306.5,-168.5</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1063</ID>
<type>DA_FROM</type>
<position>497.5,-60</position>
<input>
<ID>IN_0</ID>1056 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>285</ID>
<type>DA_FROM</type>
<position>306.5,-171.5</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1064</ID>
<type>DA_FROM</type>
<position>497.5,-63</position>
<input>
<ID>IN_0</ID>1057 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>286</ID>
<type>DA_FROM</type>
<position>306.5,-174</position>
<input>
<ID>IN_0</ID>257 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1065</ID>
<type>DA_FROM</type>
<position>497.5,-65.5</position>
<input>
<ID>IN_0</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>287</ID>
<type>DA_FROM</type>
<position>307,-177</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1066</ID>
<type>DA_FROM</type>
<position>498,-68.5</position>
<input>
<ID>IN_0</ID>1059 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>288</ID>
<type>DA_FROM</type>
<position>307,-179.5</position>
<input>
<ID>IN_0</ID>259 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>1067</ID>
<type>DA_FROM</type>
<position>498,-71</position>
<input>
<ID>IN_0</ID>1060 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>289</ID>
<type>DE_TO</type>
<position>335.5,-168</position>
<input>
<ID>IN_0</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BUS-PC</lparam></gate>
<gate>
<ID>1068</ID>
<type>DE_TO</type>
<position>526.5,-59.5</position>
<input>
<ID>IN_0</ID>1061 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SP-DEC</lparam></gate>
<gate>
<ID>324</ID>
<type>AA_LABEL</type>
<position>158,-39</position>
<gparam>LABEL_TEXT Conditionals</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>325</ID>
<type>DE_OR8</type>
<position>180.5,-61.5</position>
<input>
<ID>IN_0</ID>367 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>339 </input>
<input>
<ID>IN_3</ID>340 </input>
<input>
<ID>IN_4</ID>359 </input>
<input>
<ID>IN_5</ID>358 </input>
<input>
<ID>IN_6</ID>342 </input>
<input>
<ID>IN_7</ID>341 </input>
<output>
<ID>OUT</ID>360 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>326</ID>
<type>DA_FROM</type>
<position>160.5,-47.5</position>
<input>
<ID>IN_0</ID>361 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZ</lparam></gate>
<gate>
<ID>328</ID>
<type>DA_FROM</type>
<position>161,-59.5</position>
<input>
<ID>IN_0</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>329</ID>
<type>DA_FROM</type>
<position>161,-62</position>
<input>
<ID>IN_0</ID>340 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>330</ID>
<type>DA_FROM</type>
<position>161,-65</position>
<input>
<ID>IN_0</ID>341 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>331</ID>
<type>DA_FROM</type>
<position>161,-67.5</position>
<input>
<ID>IN_0</ID>342 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>332</ID>
<type>DA_FROM</type>
<position>161.5,-70.5</position>
<input>
<ID>IN_0</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>333</ID>
<type>DA_FROM</type>
<position>161.5,-73</position>
<input>
<ID>IN_0</ID>359 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>334</ID>
<type>DE_TO</type>
<position>190,-61.5</position>
<input>
<ID>IN_0</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BRA</lparam></gate>
<gate>
<ID>726</ID>
<type>DE_OR8</type>
<position>327,-198</position>
<input>
<ID>IN_0</ID>730 </input>
<input>
<ID>IN_1</ID>731 </input>
<input>
<ID>IN_2</ID>732 </input>
<input>
<ID>IN_3</ID>733 </input>
<input>
<ID>IN_4</ID>737 </input>
<input>
<ID>IN_5</ID>736 </input>
<input>
<ID>IN_6</ID>735 </input>
<input>
<ID>IN_7</ID>734 </input>
<output>
<ID>OUT</ID>738 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>728</ID>
<type>DA_FROM</type>
<position>317,-191</position>
<input>
<ID>IN_0</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>730</ID>
<type>DA_FROM</type>
<position>309,-193.5</position>
<input>
<ID>IN_0</ID>731 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>731</ID>
<type>DA_FROM</type>
<position>307.5,-196</position>
<input>
<ID>IN_0</ID>732 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>732</ID>
<type>DA_FROM</type>
<position>307.5,-198.5</position>
<input>
<ID>IN_0</ID>733 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>733</ID>
<type>DA_FROM</type>
<position>307.5,-201.5</position>
<input>
<ID>IN_0</ID>734 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>738</ID>
<type>DA_FROM</type>
<position>307.5,-204</position>
<input>
<ID>IN_0</ID>735 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>742</ID>
<type>DA_FROM</type>
<position>308,-207</position>
<input>
<ID>IN_0</ID>736 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>743</ID>
<type>DA_FROM</type>
<position>308,-209.5</position>
<input>
<ID>IN_0</ID>737 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>744</ID>
<type>DE_TO</type>
<position>336.5,-198</position>
<input>
<ID>IN_0</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-ADDR</lparam></gate>
<gate>
<ID>361</ID>
<type>DA_FROM</type>
<position>153.5,-51.5</position>
<input>
<ID>IN_0</ID>366 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Zero</lparam></gate>
<gate>
<ID>365</ID>
<type>AA_AND2</type>
<position>168.5,-50</position>
<input>
<ID>IN_0</ID>361 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>367 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-59,171,-56</points>
<intersection>-59 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-56,171,-56</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>171 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>171,-59,177.5,-59</points>
<connection>
<GID>325</GID>
<name>IN_1</name></connection>
<intersection>171 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162.5,-55,163.5,-55</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>816</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>384.5,-121,389.5,-121</points>
<connection>
<GID>831</GID>
<name>IN_0</name></connection>
<intersection>389.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>389.5,-124.5,389.5,-121</points>
<connection>
<GID>830</GID>
<name>IN_0</name></connection>
<intersection>-121 1</intersection></vsegment></shape></wire>
<wire>
<ID>817</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>376.5,-123.5,388,-123.5</points>
<connection>
<GID>832</GID>
<name>IN_0</name></connection>
<intersection>388 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>388,-125.5,388,-123.5</points>
<intersection>-125.5 8</intersection>
<intersection>-123.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>388,-125.5,389.5,-125.5</points>
<connection>
<GID>830</GID>
<name>IN_1</name></connection>
<intersection>388 7</intersection></hsegment></shape></wire>
<wire>
<ID>818</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>387,-126.5,387,-126</points>
<intersection>-126.5 1</intersection>
<intersection>-126 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>387,-126.5,389.5,-126.5</points>
<connection>
<GID>830</GID>
<name>IN_2</name></connection>
<intersection>387 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375,-126,387,-126</points>
<connection>
<GID>833</GID>
<name>IN_0</name></connection>
<intersection>387 0</intersection></hsegment></shape></wire>
<wire>
<ID>819</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>377,-128.5,377,-127.5</points>
<intersection>-128.5 2</intersection>
<intersection>-127.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>377,-127.5,389.5,-127.5</points>
<connection>
<GID>830</GID>
<name>IN_3</name></connection>
<intersection>377 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375,-128.5,377,-128.5</points>
<connection>
<GID>834</GID>
<name>IN_0</name></connection>
<intersection>377 0</intersection></hsegment></shape></wire>
<wire>
<ID>820</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>378,-131.5,378,-128.5</points>
<intersection>-131.5 2</intersection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>378,-128.5,389.5,-128.5</points>
<connection>
<GID>830</GID>
<name>IN_7</name></connection>
<intersection>378 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375,-131.5,378,-131.5</points>
<connection>
<GID>835</GID>
<name>IN_0</name></connection>
<intersection>378 0</intersection></hsegment></shape></wire>
<wire>
<ID>821</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379.5,-134,379.5,-129.5</points>
<intersection>-134 2</intersection>
<intersection>-129.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379.5,-129.5,389.5,-129.5</points>
<connection>
<GID>830</GID>
<name>IN_6</name></connection>
<intersection>379.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375,-134,379.5,-134</points>
<connection>
<GID>836</GID>
<name>IN_0</name></connection>
<intersection>379.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>822</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381.5,-137,381.5,-130.5</points>
<intersection>-137 2</intersection>
<intersection>-130.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381.5,-130.5,389.5,-130.5</points>
<connection>
<GID>830</GID>
<name>IN_5</name></connection>
<intersection>381.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-137,381.5,-137</points>
<connection>
<GID>837</GID>
<name>IN_0</name></connection>
<intersection>381.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>823</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>383.5,-139.5,383.5,-131.5</points>
<intersection>-139.5 2</intersection>
<intersection>-131.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>383.5,-131.5,389.5,-131.5</points>
<connection>
<GID>830</GID>
<name>IN_4</name></connection>
<intersection>383.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-139.5,383.5,-139.5</points>
<connection>
<GID>838</GID>
<name>IN_0</name></connection>
<intersection>383.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>824</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>396.5,-128,400,-128</points>
<connection>
<GID>830</GID>
<name>OUT</name></connection>
<connection>
<GID>839</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>825</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382,-55,387,-55</points>
<connection>
<GID>841</GID>
<name>IN_0</name></connection>
<intersection>387 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>387,-58.5,387,-55</points>
<connection>
<GID>840</GID>
<name>IN_0</name></connection>
<intersection>-55 1</intersection></vsegment></shape></wire>
<wire>
<ID>826</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>374,-57.5,385.5,-57.5</points>
<connection>
<GID>842</GID>
<name>IN_0</name></connection>
<intersection>385.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>385.5,-59.5,385.5,-57.5</points>
<intersection>-59.5 8</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>385.5,-59.5,387,-59.5</points>
<connection>
<GID>840</GID>
<name>IN_1</name></connection>
<intersection>385.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>827</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384.5,-60.5,384.5,-60</points>
<intersection>-60.5 1</intersection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384.5,-60.5,387,-60.5</points>
<connection>
<GID>840</GID>
<name>IN_2</name></connection>
<intersection>384.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-60,384.5,-60</points>
<connection>
<GID>843</GID>
<name>IN_0</name></connection>
<intersection>384.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>828</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374.5,-62.5,374.5,-61.5</points>
<intersection>-62.5 2</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>374.5,-61.5,387,-61.5</points>
<connection>
<GID>840</GID>
<name>IN_3</name></connection>
<intersection>374.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-62.5,374.5,-62.5</points>
<connection>
<GID>844</GID>
<name>IN_0</name></connection>
<intersection>374.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>829</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375.5,-65.5,375.5,-62.5</points>
<intersection>-65.5 2</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375.5,-62.5,387,-62.5</points>
<connection>
<GID>840</GID>
<name>IN_7</name></connection>
<intersection>375.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-65.5,375.5,-65.5</points>
<connection>
<GID>845</GID>
<name>IN_0</name></connection>
<intersection>375.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>830</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>377,-68,377,-63.5</points>
<intersection>-68 2</intersection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>377,-63.5,387,-63.5</points>
<connection>
<GID>840</GID>
<name>IN_6</name></connection>
<intersection>377 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-68,377,-68</points>
<connection>
<GID>846</GID>
<name>IN_0</name></connection>
<intersection>377 0</intersection></hsegment></shape></wire>
<wire>
<ID>831</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379,-71,379,-64.5</points>
<intersection>-71 2</intersection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,-64.5,387,-64.5</points>
<connection>
<GID>840</GID>
<name>IN_5</name></connection>
<intersection>379 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>373,-71,379,-71</points>
<connection>
<GID>847</GID>
<name>IN_0</name></connection>
<intersection>379 0</intersection></hsegment></shape></wire>
<wire>
<ID>832</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381,-73.5,381,-65.5</points>
<intersection>-73.5 2</intersection>
<intersection>-65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381,-65.5,387,-65.5</points>
<connection>
<GID>840</GID>
<name>IN_4</name></connection>
<intersection>381 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>373,-73.5,381,-73.5</points>
<connection>
<GID>848</GID>
<name>IN_0</name></connection>
<intersection>381 0</intersection></hsegment></shape></wire>
<wire>
<ID>833</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>394,-62,397.5,-62</points>
<connection>
<GID>840</GID>
<name>OUT</name></connection>
<connection>
<GID>849</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>834</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382,-86.5,387,-86.5</points>
<connection>
<GID>851</GID>
<name>IN_0</name></connection>
<intersection>387 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>387,-90,387,-86.5</points>
<connection>
<GID>850</GID>
<name>IN_0</name></connection>
<intersection>-86.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>835</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>374,-89,385.5,-89</points>
<connection>
<GID>852</GID>
<name>IN_0</name></connection>
<intersection>385.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>385.5,-91,385.5,-89</points>
<intersection>-91 8</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>385.5,-91,387,-91</points>
<connection>
<GID>850</GID>
<name>IN_1</name></connection>
<intersection>385.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>836</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384.5,-92,384.5,-91.5</points>
<intersection>-92 1</intersection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384.5,-92,387,-92</points>
<connection>
<GID>850</GID>
<name>IN_2</name></connection>
<intersection>384.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-91.5,384.5,-91.5</points>
<connection>
<GID>853</GID>
<name>IN_0</name></connection>
<intersection>384.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>837</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374.5,-94,374.5,-93</points>
<intersection>-94 2</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>374.5,-93,387,-93</points>
<connection>
<GID>850</GID>
<name>IN_3</name></connection>
<intersection>374.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-94,374.5,-94</points>
<connection>
<GID>854</GID>
<name>IN_0</name></connection>
<intersection>374.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>838</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375.5,-97,375.5,-94</points>
<intersection>-97 2</intersection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375.5,-94,387,-94</points>
<connection>
<GID>850</GID>
<name>IN_7</name></connection>
<intersection>375.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-97,375.5,-97</points>
<connection>
<GID>855</GID>
<name>IN_0</name></connection>
<intersection>375.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>839</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>377,-99.5,377,-95</points>
<intersection>-99.5 2</intersection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>377,-95,387,-95</points>
<connection>
<GID>850</GID>
<name>IN_6</name></connection>
<intersection>377 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-99.5,377,-99.5</points>
<connection>
<GID>856</GID>
<name>IN_0</name></connection>
<intersection>377 0</intersection></hsegment></shape></wire>
<wire>
<ID>840</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379,-102.5,379,-96</points>
<intersection>-102.5 2</intersection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,-96,387,-96</points>
<connection>
<GID>850</GID>
<name>IN_5</name></connection>
<intersection>379 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>373,-102.5,379,-102.5</points>
<connection>
<GID>857</GID>
<name>IN_0</name></connection>
<intersection>379 0</intersection></hsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-248.5,129,-248.5</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>129 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>129,-252,129,-248.5</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>-248.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>841</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381,-105,381,-97</points>
<intersection>-105 2</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381,-97,387,-97</points>
<connection>
<GID>850</GID>
<name>IN_4</name></connection>
<intersection>381 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>373,-105,381,-105</points>
<connection>
<GID>858</GID>
<name>IN_0</name></connection>
<intersection>381 0</intersection></hsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,-251,127.5,-251</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>127.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>127.5,-253,127.5,-251</points>
<intersection>-253 8</intersection>
<intersection>-251 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>127.5,-253,129,-253</points>
<connection>
<GID>414</GID>
<name>IN_1</name></connection>
<intersection>127.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>842</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>394,-93.5,397.5,-93.5</points>
<connection>
<GID>850</GID>
<name>OUT</name></connection>
<connection>
<GID>859</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-254,126.5,-253.5</points>
<intersection>-254 1</intersection>
<intersection>-253.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126.5,-254,129,-254</points>
<connection>
<GID>414</GID>
<name>IN_2</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-253.5,126.5,-253.5</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>843</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>385,-152.5,390,-152.5</points>
<connection>
<GID>861</GID>
<name>IN_0</name></connection>
<intersection>390 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>390,-156,390,-152.5</points>
<connection>
<GID>860</GID>
<name>IN_0</name></connection>
<intersection>-152.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-256,116.5,-255</points>
<intersection>-256 2</intersection>
<intersection>-255 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-255,129,-255</points>
<connection>
<GID>414</GID>
<name>IN_3</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-256,116.5,-256</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>844</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>377,-155,388.5,-155</points>
<connection>
<GID>862</GID>
<name>IN_0</name></connection>
<intersection>388.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>388.5,-157,388.5,-155</points>
<intersection>-157 8</intersection>
<intersection>-155 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>388.5,-157,390,-157</points>
<connection>
<GID>860</GID>
<name>IN_1</name></connection>
<intersection>388.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>845</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>387.5,-158,387.5,-157.5</points>
<intersection>-158 1</intersection>
<intersection>-157.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>387.5,-158,390,-158</points>
<connection>
<GID>860</GID>
<name>IN_2</name></connection>
<intersection>387.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-157.5,387.5,-157.5</points>
<connection>
<GID>863</GID>
<name>IN_0</name></connection>
<intersection>387.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>846</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>377.5,-160,377.5,-159</points>
<intersection>-160 2</intersection>
<intersection>-159 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>377.5,-159,390,-159</points>
<connection>
<GID>860</GID>
<name>IN_3</name></connection>
<intersection>377.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-160,377.5,-160</points>
<connection>
<GID>864</GID>
<name>IN_0</name></connection>
<intersection>377.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>847</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>378.5,-163,378.5,-160</points>
<intersection>-163 2</intersection>
<intersection>-160 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>378.5,-160,390,-160</points>
<connection>
<GID>860</GID>
<name>IN_7</name></connection>
<intersection>378.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-163,378.5,-163</points>
<connection>
<GID>865</GID>
<name>IN_0</name></connection>
<intersection>378.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>848</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380,-165.5,380,-161</points>
<intersection>-165.5 2</intersection>
<intersection>-161 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380,-161,390,-161</points>
<connection>
<GID>860</GID>
<name>IN_6</name></connection>
<intersection>380 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-165.5,380,-165.5</points>
<connection>
<GID>866</GID>
<name>IN_0</name></connection>
<intersection>380 0</intersection></hsegment></shape></wire>
<wire>
<ID>849</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>382,-168.5,382,-162</points>
<intersection>-168.5 2</intersection>
<intersection>-162 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>382,-162,390,-162</points>
<connection>
<GID>860</GID>
<name>IN_5</name></connection>
<intersection>382 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>376,-168.5,382,-168.5</points>
<connection>
<GID>867</GID>
<name>IN_0</name></connection>
<intersection>382 0</intersection></hsegment></shape></wire>
<wire>
<ID>850</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384,-171,384,-163</points>
<intersection>-171 2</intersection>
<intersection>-163 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384,-163,390,-163</points>
<connection>
<GID>860</GID>
<name>IN_4</name></connection>
<intersection>384 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>376,-171,384,-171</points>
<connection>
<GID>868</GID>
<name>IN_0</name></connection>
<intersection>384 0</intersection></hsegment></shape></wire>
<wire>
<ID>851</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>397,-159.5,400.5,-159.5</points>
<connection>
<GID>869</GID>
<name>IN_0</name></connection>
<connection>
<GID>860</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>852</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>385,-178.5,390,-178.5</points>
<connection>
<GID>876</GID>
<name>IN_0</name></connection>
<intersection>390 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>390,-182,390,-178.5</points>
<connection>
<GID>875</GID>
<name>IN_0</name></connection>
<intersection>-178.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>853</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>377,-181,388.5,-181</points>
<connection>
<GID>877</GID>
<name>IN_0</name></connection>
<intersection>388.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>388.5,-183,388.5,-181</points>
<intersection>-183 8</intersection>
<intersection>-181 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>388.5,-183,390,-183</points>
<connection>
<GID>875</GID>
<name>IN_1</name></connection>
<intersection>388.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>854</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>387.5,-184,387.5,-183.5</points>
<intersection>-184 1</intersection>
<intersection>-183.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>387.5,-184,390,-184</points>
<connection>
<GID>875</GID>
<name>IN_2</name></connection>
<intersection>387.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-183.5,387.5,-183.5</points>
<connection>
<GID>878</GID>
<name>IN_0</name></connection>
<intersection>387.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>855</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>377.5,-186,377.5,-185</points>
<intersection>-186 2</intersection>
<intersection>-185 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>377.5,-185,390,-185</points>
<connection>
<GID>875</GID>
<name>IN_3</name></connection>
<intersection>377.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-186,377.5,-186</points>
<connection>
<GID>879</GID>
<name>IN_0</name></connection>
<intersection>377.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>856</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>378.5,-189,378.5,-186</points>
<intersection>-189 2</intersection>
<intersection>-186 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>378.5,-186,390,-186</points>
<connection>
<GID>875</GID>
<name>IN_7</name></connection>
<intersection>378.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-189,378.5,-189</points>
<connection>
<GID>880</GID>
<name>IN_0</name></connection>
<intersection>378.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>857</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380,-191.5,380,-187</points>
<intersection>-191.5 2</intersection>
<intersection>-187 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380,-187,390,-187</points>
<connection>
<GID>875</GID>
<name>IN_6</name></connection>
<intersection>380 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-191.5,380,-191.5</points>
<connection>
<GID>881</GID>
<name>IN_0</name></connection>
<intersection>380 0</intersection></hsegment></shape></wire>
<wire>
<ID>858</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>382,-194.5,382,-188</points>
<intersection>-194.5 2</intersection>
<intersection>-188 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>382,-188,390,-188</points>
<connection>
<GID>875</GID>
<name>IN_5</name></connection>
<intersection>382 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>376,-194.5,382,-194.5</points>
<connection>
<GID>882</GID>
<name>IN_0</name></connection>
<intersection>382 0</intersection></hsegment></shape></wire>
<wire>
<ID>859</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384,-197,384,-189</points>
<intersection>-197 2</intersection>
<intersection>-189 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384,-189,390,-189</points>
<connection>
<GID>875</GID>
<name>IN_4</name></connection>
<intersection>384 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>376,-197,384,-197</points>
<connection>
<GID>883</GID>
<name>IN_0</name></connection>
<intersection>384 0</intersection></hsegment></shape></wire>
<wire>
<ID>860</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>397,-185.5,400.5,-185.5</points>
<connection>
<GID>875</GID>
<name>OUT</name></connection>
<connection>
<GID>884</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>861</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382,-208.5,387,-208.5</points>
<connection>
<GID>887</GID>
<name>IN_0</name></connection>
<intersection>387 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>387,-212,387,-208.5</points>
<connection>
<GID>886</GID>
<name>IN_0</name></connection>
<intersection>-208.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>862</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>374,-211,385.5,-211</points>
<connection>
<GID>888</GID>
<name>IN_0</name></connection>
<intersection>385.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>385.5,-213,385.5,-211</points>
<intersection>-213 8</intersection>
<intersection>-211 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>385.5,-213,387,-213</points>
<connection>
<GID>886</GID>
<name>IN_1</name></connection>
<intersection>385.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>863</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384.5,-214,384.5,-213.5</points>
<intersection>-214 1</intersection>
<intersection>-213.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384.5,-214,387,-214</points>
<connection>
<GID>886</GID>
<name>IN_2</name></connection>
<intersection>384.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-213.5,384.5,-213.5</points>
<connection>
<GID>889</GID>
<name>IN_0</name></connection>
<intersection>384.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>864</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374.5,-216,374.5,-215</points>
<intersection>-216 2</intersection>
<intersection>-215 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>374.5,-215,387,-215</points>
<connection>
<GID>886</GID>
<name>IN_3</name></connection>
<intersection>374.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-216,374.5,-216</points>
<connection>
<GID>890</GID>
<name>IN_0</name></connection>
<intersection>374.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>865</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375.5,-219,375.5,-216</points>
<intersection>-219 2</intersection>
<intersection>-216 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375.5,-216,387,-216</points>
<connection>
<GID>886</GID>
<name>IN_7</name></connection>
<intersection>375.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-219,375.5,-219</points>
<connection>
<GID>891</GID>
<name>IN_0</name></connection>
<intersection>375.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>866</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>377,-221.5,377,-217</points>
<intersection>-221.5 2</intersection>
<intersection>-217 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>377,-217,387,-217</points>
<connection>
<GID>886</GID>
<name>IN_6</name></connection>
<intersection>377 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-221.5,377,-221.5</points>
<connection>
<GID>892</GID>
<name>IN_0</name></connection>
<intersection>377 0</intersection></hsegment></shape></wire>
<wire>
<ID>867</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379,-224.5,379,-218</points>
<intersection>-224.5 2</intersection>
<intersection>-218 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379,-218,387,-218</points>
<connection>
<GID>886</GID>
<name>IN_5</name></connection>
<intersection>379 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>373,-224.5,379,-224.5</points>
<connection>
<GID>893</GID>
<name>IN_0</name></connection>
<intersection>379 0</intersection></hsegment></shape></wire>
<wire>
<ID>868</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381,-227,381,-219</points>
<intersection>-227 2</intersection>
<intersection>-219 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381,-219,387,-219</points>
<connection>
<GID>886</GID>
<name>IN_4</name></connection>
<intersection>381 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>373,-227,381,-227</points>
<connection>
<GID>894</GID>
<name>IN_0</name></connection>
<intersection>381 0</intersection></hsegment></shape></wire>
<wire>
<ID>869</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>394,-215.5,397.5,-215.5</points>
<connection>
<GID>886</GID>
<name>OUT</name></connection>
<connection>
<GID>895</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>871</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>451.5,-121,463,-121</points>
<connection>
<GID>961</GID>
<name>IN_0</name></connection>
<intersection>463 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>463,-123,463,-121</points>
<intersection>-123 8</intersection>
<intersection>-121 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>463,-123,464.5,-123</points>
<connection>
<GID>900</GID>
<name>IN_1</name></connection>
<intersection>463 7</intersection></hsegment></shape></wire>
<wire>
<ID>872</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462,-124,462,-123.5</points>
<intersection>-124 1</intersection>
<intersection>-123.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>462,-124,464.5,-124</points>
<connection>
<GID>900</GID>
<name>IN_2</name></connection>
<intersection>462 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450,-123.5,462,-123.5</points>
<connection>
<GID>969</GID>
<name>IN_0</name></connection>
<intersection>462 0</intersection></hsegment></shape></wire>
<wire>
<ID>873</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452,-126,452,-125</points>
<intersection>-126 2</intersection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>452,-125,464.5,-125</points>
<connection>
<GID>900</GID>
<name>IN_3</name></connection>
<intersection>452 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450,-126,452,-126</points>
<connection>
<GID>981</GID>
<name>IN_0</name></connection>
<intersection>452 0</intersection></hsegment></shape></wire>
<wire>
<ID>874</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>453,-129,453,-126</points>
<intersection>-129 2</intersection>
<intersection>-126 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>453,-126,464.5,-126</points>
<connection>
<GID>900</GID>
<name>IN_7</name></connection>
<intersection>453 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450,-129,453,-129</points>
<connection>
<GID>982</GID>
<name>IN_0</name></connection>
<intersection>453 0</intersection></hsegment></shape></wire>
<wire>
<ID>875</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454.5,-131.5,454.5,-127</points>
<intersection>-131.5 2</intersection>
<intersection>-127 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>454.5,-127,464.5,-127</points>
<connection>
<GID>900</GID>
<name>IN_6</name></connection>
<intersection>454.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450,-131.5,454.5,-131.5</points>
<connection>
<GID>983</GID>
<name>IN_0</name></connection>
<intersection>454.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>876</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456.5,-134.5,456.5,-128</points>
<intersection>-134.5 2</intersection>
<intersection>-128 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>456.5,-128,464.5,-128</points>
<connection>
<GID>900</GID>
<name>IN_5</name></connection>
<intersection>456.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450.5,-134.5,456.5,-134.5</points>
<connection>
<GID>985</GID>
<name>IN_0</name></connection>
<intersection>456.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>877</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458.5,-137,458.5,-129</points>
<intersection>-137 2</intersection>
<intersection>-129 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>458.5,-129,464.5,-129</points>
<connection>
<GID>900</GID>
<name>IN_4</name></connection>
<intersection>458.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450.5,-137,458.5,-137</points>
<connection>
<GID>987</GID>
<name>IN_0</name></connection>
<intersection>458.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>878</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>471.5,-125.5,475,-125.5</points>
<connection>
<GID>900</GID>
<name>OUT</name></connection>
<connection>
<GID>989</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-259,117.5,-256</points>
<intersection>-259 2</intersection>
<intersection>-256 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-256,129,-256</points>
<connection>
<GID>414</GID>
<name>IN_7</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-259,117.5,-259</points>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-261.5,119,-257</points>
<intersection>-261.5 2</intersection>
<intersection>-257 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-257,129,-257</points>
<connection>
<GID>414</GID>
<name>IN_6</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-261.5,119,-261.5</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-264.5,121,-258</points>
<intersection>-264.5 2</intersection>
<intersection>-258 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-258,129,-258</points>
<connection>
<GID>414</GID>
<name>IN_5</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-264.5,121,-264.5</points>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-267,123,-259</points>
<intersection>-267 2</intersection>
<intersection>-259 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-259,129,-259</points>
<connection>
<GID>414</GID>
<name>IN_4</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-267,123,-267</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>902</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>457,-52.5,462,-52.5</points>
<connection>
<GID>993</GID>
<name>IN_0</name></connection>
<intersection>462 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>462,-56,462,-52.5</points>
<connection>
<GID>991</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>905</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>381.5,-233,386.5,-233</points>
<connection>
<GID>936</GID>
<name>IN_0</name></connection>
<intersection>386.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>386.5,-236.5,386.5,-233</points>
<connection>
<GID>935</GID>
<name>IN_0</name></connection>
<intersection>-233 1</intersection></vsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>155.5,-57,163.5,-57</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<connection>
<GID>56</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>906</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>373.5,-235.5,385,-235.5</points>
<connection>
<GID>937</GID>
<name>IN_0</name></connection>
<intersection>385 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>385,-237.5,385,-235.5</points>
<intersection>-237.5 8</intersection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>385,-237.5,386.5,-237.5</points>
<connection>
<GID>935</GID>
<name>IN_1</name></connection>
<intersection>385 7</intersection></hsegment></shape></wire>
<wire>
<ID>907</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384,-238.5,384,-238</points>
<intersection>-238.5 1</intersection>
<intersection>-238 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384,-238.5,386.5,-238.5</points>
<connection>
<GID>935</GID>
<name>IN_2</name></connection>
<intersection>384 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372,-238,384,-238</points>
<connection>
<GID>938</GID>
<name>IN_0</name></connection>
<intersection>384 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-56.5,128,-56.5</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>128 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128,-60,128,-56.5</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>-56.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>908</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374,-240.5,374,-239.5</points>
<intersection>-240.5 2</intersection>
<intersection>-239.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>374,-239.5,386.5,-239.5</points>
<connection>
<GID>935</GID>
<name>IN_3</name></connection>
<intersection>374 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372,-240.5,374,-240.5</points>
<connection>
<GID>939</GID>
<name>IN_0</name></connection>
<intersection>374 0</intersection></hsegment></shape></wire>
<wire>
<ID>909</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375,-243.5,375,-240.5</points>
<intersection>-243.5 2</intersection>
<intersection>-240.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375,-240.5,386.5,-240.5</points>
<connection>
<GID>935</GID>
<name>IN_7</name></connection>
<intersection>375 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372,-243.5,375,-243.5</points>
<connection>
<GID>940</GID>
<name>IN_0</name></connection>
<intersection>375 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115,-59,126.5,-59</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>126.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>126.5,-61,126.5,-59</points>
<intersection>-61 8</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>126.5,-61,128,-61</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>126.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>910</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>376.5,-246,376.5,-241.5</points>
<intersection>-246 2</intersection>
<intersection>-241.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>376.5,-241.5,386.5,-241.5</points>
<connection>
<GID>935</GID>
<name>IN_6</name></connection>
<intersection>376.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372,-246,376.5,-246</points>
<connection>
<GID>941</GID>
<name>IN_0</name></connection>
<intersection>376.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-3,32,-3</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>911</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>378.5,-249,378.5,-242.5</points>
<intersection>-249 2</intersection>
<intersection>-242.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>378.5,-242.5,386.5,-242.5</points>
<connection>
<GID>935</GID>
<name>IN_5</name></connection>
<intersection>378.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-249,378.5,-249</points>
<connection>
<GID>942</GID>
<name>IN_0</name></connection>
<intersection>378.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-62,125.5,-61.5</points>
<intersection>-62 1</intersection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125.5,-62,128,-62</points>
<connection>
<GID>152</GID>
<name>IN_2</name></connection>
<intersection>125.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-61.5,125.5,-61.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>912</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380.5,-251.5,380.5,-243.5</points>
<intersection>-251.5 2</intersection>
<intersection>-243.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380.5,-243.5,386.5,-243.5</points>
<connection>
<GID>935</GID>
<name>IN_4</name></connection>
<intersection>380.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>372.5,-251.5,380.5,-251.5</points>
<connection>
<GID>943</GID>
<name>IN_0</name></connection>
<intersection>380.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-64,115.5,-63</points>
<intersection>-64 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-63,128,-63</points>
<connection>
<GID>152</GID>
<name>IN_3</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-64,115.5,-64</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>913</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>393.5,-240,397,-240</points>
<connection>
<GID>944</GID>
<name>IN_0</name></connection>
<connection>
<GID>935</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-67,116.5,-64</points>
<intersection>-67 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-64,128,-64</points>
<connection>
<GID>152</GID>
<name>IN_7</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-67,116.5,-67</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>914</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>449,-55,460.5,-55</points>
<connection>
<GID>995</GID>
<name>IN_0</name></connection>
<intersection>460.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>460.5,-57,460.5,-55</points>
<intersection>-57 8</intersection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>460.5,-57,462,-57</points>
<connection>
<GID>991</GID>
<name>IN_1</name></connection>
<intersection>460.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>136,-255.5,139.5,-255.5</points>
<connection>
<GID>414</GID>
<name>OUT</name></connection>
<connection>
<GID>460</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-69.5,118,-65</points>
<intersection>-69.5 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-65,128,-65</points>
<connection>
<GID>152</GID>
<name>IN_6</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-69.5,118,-69.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>915</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459.5,-58,459.5,-57.5</points>
<intersection>-58 1</intersection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>459.5,-58,462,-58</points>
<connection>
<GID>991</GID>
<name>IN_2</name></connection>
<intersection>459.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-57.5,459.5,-57.5</points>
<connection>
<GID>997</GID>
<name>IN_0</name></connection>
<intersection>459.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-214,129,-214</points>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<intersection>129 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>129,-217.5,129,-214</points>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<intersection>-214 1</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-72.5,120,-66</points>
<intersection>-72.5 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-66,128,-66</points>
<connection>
<GID>152</GID>
<name>IN_5</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-72.5,120,-72.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>916</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449.5,-60,449.5,-59</points>
<intersection>-60 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>449.5,-59,462,-59</points>
<connection>
<GID>991</GID>
<name>IN_3</name></connection>
<intersection>449.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-60,449.5,-60</points>
<connection>
<GID>1000</GID>
<name>IN_0</name></connection>
<intersection>449.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,-216.5,127.5,-216.5</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>127.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>127.5,-218.5,127.5,-216.5</points>
<intersection>-218.5 8</intersection>
<intersection>-216.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>127.5,-218.5,129,-218.5</points>
<connection>
<GID>445</GID>
<name>IN_1</name></connection>
<intersection>127.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-75,122,-67</points>
<intersection>-75 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,-67,128,-67</points>
<connection>
<GID>152</GID>
<name>IN_4</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-75,122,-75</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>917</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>450.5,-63,450.5,-60</points>
<intersection>-63 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>450.5,-60,462,-60</points>
<connection>
<GID>991</GID>
<name>IN_7</name></connection>
<intersection>450.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-63,450.5,-63</points>
<connection>
<GID>1002</GID>
<name>IN_0</name></connection>
<intersection>450.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-219.5,126.5,-219</points>
<intersection>-219.5 1</intersection>
<intersection>-219 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126.5,-219.5,129,-219.5</points>
<connection>
<GID>445</GID>
<name>IN_2</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-219,126.5,-219</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135,-63.5,138.5,-63.5</points>
<connection>
<GID>152</GID>
<name>OUT</name></connection>
<connection>
<GID>169</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-221.5,116.5,-220.5</points>
<intersection>-221.5 2</intersection>
<intersection>-220.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-220.5,129,-220.5</points>
<connection>
<GID>445</GID>
<name>IN_3</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-221.5,116.5,-221.5</points>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-84.5,129,-84.5</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>129 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>129,-88,129,-84.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>-84.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-224.5,117.5,-221.5</points>
<intersection>-224.5 2</intersection>
<intersection>-221.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-221.5,129,-221.5</points>
<connection>
<GID>445</GID>
<name>IN_7</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-224.5,117.5,-224.5</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,-87,127.5,-87</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>127.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>127.5,-89,127.5,-87</points>
<intersection>-89 8</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>127.5,-89,129,-89</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>127.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-90,126.5,-89.5</points>
<intersection>-90 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126.5,-90,129,-90</points>
<connection>
<GID>170</GID>
<name>IN_2</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-89.5,126.5,-89.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-92,116.5,-91</points>
<intersection>-92 2</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-91,129,-91</points>
<connection>
<GID>170</GID>
<name>IN_3</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-92,116.5,-92</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-95,117.5,-92</points>
<intersection>-95 2</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-92,129,-92</points>
<connection>
<GID>170</GID>
<name>IN_7</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-95,117.5,-95</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-97.5,119,-93</points>
<intersection>-97.5 2</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-93,129,-93</points>
<connection>
<GID>170</GID>
<name>IN_6</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-97.5,119,-97.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-100.5,121,-94</points>
<intersection>-100.5 2</intersection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-94,129,-94</points>
<connection>
<GID>170</GID>
<name>IN_5</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-100.5,121,-100.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-103,123,-95</points>
<intersection>-103 2</intersection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-95,129,-95</points>
<connection>
<GID>170</GID>
<name>IN_4</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-103,123,-103</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>136,-91.5,139.5,-91.5</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<connection>
<GID>179</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225.5,-122.5,230.5,-122.5</points>
<connection>
<GID>611</GID>
<name>IN_0</name></connection>
<intersection>230.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>230.5,-126,230.5,-122.5</points>
<connection>
<GID>610</GID>
<name>IN_0</name></connection>
<intersection>-122.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-129,30.5,-129</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>30.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>30.5,-132.5,30.5,-129</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>-129 1</intersection></vsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217.5,-125,229,-125</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>229 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>229,-127,229,-125</points>
<intersection>-127 8</intersection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>229,-127,230.5,-127</points>
<connection>
<GID>610</GID>
<name>IN_1</name></connection>
<intersection>229 7</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-131.5,29,-131.5</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>29 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>29,-133.5,29,-131.5</points>
<intersection>-133.5 8</intersection>
<intersection>-131.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>29,-133.5,30.5,-133.5</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>29 7</intersection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,-128,228,-127.5</points>
<intersection>-128 1</intersection>
<intersection>-127.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>228,-128,230.5,-128</points>
<connection>
<GID>610</GID>
<name>IN_2</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-127.5,228,-127.5</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-134.5,28,-134</points>
<intersection>-134.5 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-134.5,30.5,-134.5</points>
<connection>
<GID>180</GID>
<name>IN_2</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-134,28,-134</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-130,218,-129</points>
<intersection>-130 2</intersection>
<intersection>-129 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-129,230.5,-129</points>
<connection>
<GID>610</GID>
<name>IN_3</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-130,218,-130</points>
<connection>
<GID>614</GID>
<name>IN_0</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-136.5,18,-135.5</points>
<intersection>-136.5 2</intersection>
<intersection>-135.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-135.5,30.5,-135.5</points>
<connection>
<GID>180</GID>
<name>IN_3</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-136.5,18,-136.5</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-133,219,-130</points>
<intersection>-133 2</intersection>
<intersection>-130 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-130,230.5,-130</points>
<connection>
<GID>610</GID>
<name>IN_7</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-133,219,-133</points>
<connection>
<GID>615</GID>
<name>IN_0</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-139.5,19,-136.5</points>
<intersection>-139.5 2</intersection>
<intersection>-136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-136.5,30.5,-136.5</points>
<connection>
<GID>180</GID>
<name>IN_7</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-139.5,19,-139.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220.5,-135.5,220.5,-131</points>
<intersection>-135.5 2</intersection>
<intersection>-131 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>220.5,-131,230.5,-131</points>
<connection>
<GID>610</GID>
<name>IN_6</name></connection>
<intersection>220.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-135.5,220.5,-135.5</points>
<connection>
<GID>616</GID>
<name>IN_0</name></connection>
<intersection>220.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-142,20.5,-137.5</points>
<intersection>-142 2</intersection>
<intersection>-137.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-137.5,30.5,-137.5</points>
<connection>
<GID>180</GID>
<name>IN_6</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-142,20.5,-142</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,-138.5,222.5,-132</points>
<intersection>-138.5 2</intersection>
<intersection>-132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,-132,230.5,-132</points>
<connection>
<GID>610</GID>
<name>IN_5</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216.5,-138.5,222.5,-138.5</points>
<connection>
<GID>617</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-145,22.5,-138.5</points>
<intersection>-145 2</intersection>
<intersection>-138.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-138.5,30.5,-138.5</points>
<connection>
<GID>180</GID>
<name>IN_5</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-145,22.5,-145</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224.5,-141,224.5,-133</points>
<intersection>-141 2</intersection>
<intersection>-133 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224.5,-133,230.5,-133</points>
<connection>
<GID>610</GID>
<name>IN_4</name></connection>
<intersection>224.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216.5,-141,224.5,-141</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<intersection>224.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-147.5,24.5,-139.5</points>
<intersection>-147.5 2</intersection>
<intersection>-139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-139.5,30.5,-139.5</points>
<connection>
<GID>180</GID>
<name>IN_4</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-147.5,24.5,-147.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>237.5,-129.5,241,-129.5</points>
<connection>
<GID>610</GID>
<name>OUT</name></connection>
<connection>
<GID>619</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-136,41,-136</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<connection>
<GID>189</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>223,-56.5,228,-56.5</points>
<connection>
<GID>623</GID>
<name>IN_0</name></connection>
<intersection>228 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>228,-60,228,-56.5</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<intersection>-56.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-122.5,131,-122.5</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>131 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>131,-126,131,-122.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>-122.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215,-59,226.5,-59</points>
<connection>
<GID>624</GID>
<name>IN_0</name></connection>
<intersection>226.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>226.5,-61,226.5,-59</points>
<intersection>-61 8</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>226.5,-61,228,-61</points>
<connection>
<GID>622</GID>
<name>IN_1</name></connection>
<intersection>226.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118,-125,129.5,-125</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>129.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>129.5,-127,129.5,-125</points>
<intersection>-127 8</intersection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>129.5,-127,131,-127</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>129.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225.5,-62,225.5,-61.5</points>
<intersection>-62 1</intersection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225.5,-62,228,-62</points>
<connection>
<GID>622</GID>
<name>IN_2</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-61.5,225.5,-61.5</points>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<intersection>225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-128,128.5,-127.5</points>
<intersection>-128 1</intersection>
<intersection>-127.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128.5,-128,131,-128</points>
<connection>
<GID>190</GID>
<name>IN_2</name></connection>
<intersection>128.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-127.5,128.5,-127.5</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>128.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215.5,-64,215.5,-63</points>
<intersection>-64 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215.5,-63,228,-63</points>
<connection>
<GID>622</GID>
<name>IN_3</name></connection>
<intersection>215.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-64,215.5,-64</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>215.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-130,118.5,-129</points>
<intersection>-130 2</intersection>
<intersection>-129 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118.5,-129,131,-129</points>
<connection>
<GID>190</GID>
<name>IN_3</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-130,118.5,-130</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216.5,-67,216.5,-64</points>
<intersection>-67 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216.5,-64,228,-64</points>
<connection>
<GID>622</GID>
<name>IN_7</name></connection>
<intersection>216.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-67,216.5,-67</points>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<intersection>216.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-133,119.5,-130</points>
<intersection>-133 2</intersection>
<intersection>-130 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-130,131,-130</points>
<connection>
<GID>190</GID>
<name>IN_7</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-133,119.5,-133</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-69.5,218,-65</points>
<intersection>-69.5 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-65,228,-65</points>
<connection>
<GID>622</GID>
<name>IN_6</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-69.5,218,-69.5</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-135.5,121,-131</points>
<intersection>-135.5 2</intersection>
<intersection>-131 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-131,131,-131</points>
<connection>
<GID>190</GID>
<name>IN_6</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-135.5,121,-135.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,-72.5,220,-66</points>
<intersection>-72.5 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>220,-66,228,-66</points>
<connection>
<GID>622</GID>
<name>IN_5</name></connection>
<intersection>220 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214,-72.5,220,-72.5</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<intersection>220 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-138.5,123,-132</points>
<intersection>-138.5 2</intersection>
<intersection>-132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-132,131,-132</points>
<connection>
<GID>190</GID>
<name>IN_5</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>117,-138.5,123,-138.5</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-75,222,-67</points>
<intersection>-75 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222,-67,228,-67</points>
<connection>
<GID>622</GID>
<name>IN_4</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214,-75,222,-75</points>
<connection>
<GID>630</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-141,125,-133</points>
<intersection>-141 2</intersection>
<intersection>-133 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-133,131,-133</points>
<connection>
<GID>190</GID>
<name>IN_4</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>117,-141,125,-141</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235,-63.5,238.5,-63.5</points>
<connection>
<GID>622</GID>
<name>OUT</name></connection>
<connection>
<GID>631</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138,-129.5,141.5,-129.5</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<connection>
<GID>190</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>223,-88,228,-88</points>
<connection>
<GID>634</GID>
<name>IN_0</name></connection>
<intersection>228 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>228,-91.5,228,-88</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<intersection>-88 1</intersection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-59.5,30.5,-59.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>30.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>30.5,-63,30.5,-59.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-59.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215,-90.5,226.5,-90.5</points>
<connection>
<GID>635</GID>
<name>IN_0</name></connection>
<intersection>226.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>226.5,-92.5,226.5,-90.5</points>
<intersection>-92.5 8</intersection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>226.5,-92.5,228,-92.5</points>
<connection>
<GID>633</GID>
<name>IN_1</name></connection>
<intersection>226.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-62,29,-62</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>29 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>29,-64,29,-62</points>
<intersection>-64 8</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>29,-64,30.5,-64</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<intersection>29 7</intersection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225.5,-93.5,225.5,-93</points>
<intersection>-93.5 1</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225.5,-93.5,228,-93.5</points>
<connection>
<GID>633</GID>
<name>IN_2</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-93,225.5,-93</points>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<intersection>225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-65,28,-64.5</points>
<intersection>-65 1</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-65,30.5,-65</points>
<connection>
<GID>211</GID>
<name>IN_2</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-64.5,28,-64.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215.5,-95.5,215.5,-94.5</points>
<intersection>-95.5 2</intersection>
<intersection>-94.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215.5,-94.5,228,-94.5</points>
<connection>
<GID>633</GID>
<name>IN_3</name></connection>
<intersection>215.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-95.5,215.5,-95.5</points>
<connection>
<GID>637</GID>
<name>IN_0</name></connection>
<intersection>215.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-67,18,-66</points>
<intersection>-67 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-66,30.5,-66</points>
<connection>
<GID>211</GID>
<name>IN_3</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-67,18,-67</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216.5,-98.5,216.5,-95.5</points>
<intersection>-98.5 2</intersection>
<intersection>-95.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216.5,-95.5,228,-95.5</points>
<connection>
<GID>633</GID>
<name>IN_7</name></connection>
<intersection>216.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-98.5,216.5,-98.5</points>
<connection>
<GID>638</GID>
<name>IN_0</name></connection>
<intersection>216.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-70,19,-67</points>
<intersection>-70 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-67,30.5,-67</points>
<connection>
<GID>211</GID>
<name>IN_7</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-70,19,-70</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-101,218,-96.5</points>
<intersection>-101 2</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-96.5,228,-96.5</points>
<connection>
<GID>633</GID>
<name>IN_6</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-101,218,-101</points>
<connection>
<GID>639</GID>
<name>IN_0</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-72.5,20.5,-68</points>
<intersection>-72.5 2</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-68,30.5,-68</points>
<connection>
<GID>211</GID>
<name>IN_6</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-72.5,20.5,-72.5</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,-104,220,-97.5</points>
<intersection>-104 2</intersection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>220,-97.5,228,-97.5</points>
<connection>
<GID>633</GID>
<name>IN_5</name></connection>
<intersection>220 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214,-104,220,-104</points>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<intersection>220 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-75.5,22.5,-69</points>
<intersection>-75.5 2</intersection>
<intersection>-69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-69,30.5,-69</points>
<connection>
<GID>211</GID>
<name>IN_5</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-75.5,22.5,-75.5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-106.5,222,-98.5</points>
<intersection>-106.5 2</intersection>
<intersection>-98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222,-98.5,228,-98.5</points>
<connection>
<GID>633</GID>
<name>IN_4</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214,-106.5,222,-106.5</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-78,24.5,-70</points>
<intersection>-78 2</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-70,30.5,-70</points>
<connection>
<GID>211</GID>
<name>IN_4</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-78,24.5,-78</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235,-95,238.5,-95</points>
<connection>
<GID>633</GID>
<name>OUT</name></connection>
<connection>
<GID>642</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-66.5,41,-66.5</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<connection>
<GID>220</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-149.5,128,-149.5</points>
<connection>
<GID>644</GID>
<name>IN_0</name></connection>
<intersection>128 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128,-153,128,-149.5</points>
<connection>
<GID>643</GID>
<name>IN_0</name></connection>
<intersection>-149.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115,-152,126.5,-152</points>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<intersection>126.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>126.5,-154,126.5,-152</points>
<intersection>-154 8</intersection>
<intersection>-152 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>126.5,-154,128,-154</points>
<connection>
<GID>643</GID>
<name>IN_1</name></connection>
<intersection>126.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-155,125.5,-154.5</points>
<intersection>-155 1</intersection>
<intersection>-154.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125.5,-155,128,-155</points>
<connection>
<GID>643</GID>
<name>IN_2</name></connection>
<intersection>125.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-154.5,125.5,-154.5</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-157,115.5,-156</points>
<intersection>-157 2</intersection>
<intersection>-156 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-156,128,-156</points>
<connection>
<GID>643</GID>
<name>IN_3</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-157,115.5,-157</points>
<connection>
<GID>647</GID>
<name>IN_0</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-160,116.5,-157</points>
<intersection>-160 2</intersection>
<intersection>-157 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-157,128,-157</points>
<connection>
<GID>643</GID>
<name>IN_7</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-160,116.5,-160</points>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-162.5,118,-158</points>
<intersection>-162.5 2</intersection>
<intersection>-158 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-158,128,-158</points>
<connection>
<GID>643</GID>
<name>IN_6</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-162.5,118,-162.5</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-165.5,120,-159</points>
<intersection>-165.5 2</intersection>
<intersection>-159 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-159,128,-159</points>
<connection>
<GID>643</GID>
<name>IN_5</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-165.5,120,-165.5</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-168,122,-160</points>
<intersection>-168 2</intersection>
<intersection>-160 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,-160,128,-160</points>
<connection>
<GID>643</GID>
<name>IN_4</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-168,122,-168</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135,-156.5,138.5,-156.5</points>
<connection>
<GID>643</GID>
<name>OUT</name></connection>
<connection>
<GID>652</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>574</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-227,119,-222.5</points>
<intersection>-227 2</intersection>
<intersection>-222.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-222.5,129,-222.5</points>
<connection>
<GID>445</GID>
<name>IN_6</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-227,119,-227</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-230,121,-223.5</points>
<intersection>-230 2</intersection>
<intersection>-223.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-223.5,129,-223.5</points>
<connection>
<GID>445</GID>
<name>IN_5</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-230,121,-230</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-232.5,123,-224.5</points>
<intersection>-232.5 2</intersection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-224.5,129,-224.5</points>
<connection>
<GID>445</GID>
<name>IN_4</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-232.5,123,-232.5</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>136,-221,139.5,-221</points>
<connection>
<GID>445</GID>
<name>OUT</name></connection>
<connection>
<GID>470</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-92.5,30.5,-92.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>30.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>30.5,-96,30.5,-92.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-92.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-95,29,-95</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>29 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>29,-97,29,-95</points>
<intersection>-97 8</intersection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>29,-97,30.5,-97</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>29 7</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-98,28,-97.5</points>
<intersection>-98 1</intersection>
<intersection>-97.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-98,30.5,-98</points>
<connection>
<GID>118</GID>
<name>IN_2</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-97.5,28,-97.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-100,18,-99</points>
<intersection>-100 2</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-99,30.5,-99</points>
<connection>
<GID>118</GID>
<name>IN_3</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-100,18,-100</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-103,19,-100</points>
<intersection>-103 2</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-100,30.5,-100</points>
<connection>
<GID>118</GID>
<name>IN_7</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-103,19,-103</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-105.5,20.5,-101</points>
<intersection>-105.5 2</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-101,30.5,-101</points>
<connection>
<GID>118</GID>
<name>IN_6</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-105.5,20.5,-105.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-108.5,22.5,-102</points>
<intersection>-108.5 2</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-102,30.5,-102</points>
<connection>
<GID>118</GID>
<name>IN_5</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-108.5,22.5,-108.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-111,24.5,-103</points>
<intersection>-111 2</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-103,30.5,-103</points>
<connection>
<GID>118</GID>
<name>IN_4</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-111,24.5,-111</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-99.5,41,-99.5</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<connection>
<GID>149</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>317,-58,322,-58</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>322 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>322,-61.5,322,-58</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>-58 1</intersection></vsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>309,-60.5,320.5,-60.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>320.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>320.5,-62.5,320.5,-60.5</points>
<intersection>-62.5 8</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>320.5,-62.5,322,-62.5</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>320.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319.5,-63.5,319.5,-63</points>
<intersection>-63.5 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319.5,-63.5,322,-63.5</points>
<connection>
<GID>168</GID>
<name>IN_2</name></connection>
<intersection>319.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>307.5,-63,319.5,-63</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>319.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309.5,-65.5,309.5,-64.5</points>
<intersection>-65.5 2</intersection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309.5,-64.5,322,-64.5</points>
<connection>
<GID>168</GID>
<name>IN_3</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>307.5,-65.5,309.5,-65.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>309.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,-68.5,310.5,-65.5</points>
<intersection>-68.5 2</intersection>
<intersection>-65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310.5,-65.5,322,-65.5</points>
<connection>
<GID>168</GID>
<name>IN_7</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>307.5,-68.5,310.5,-68.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312,-71,312,-66.5</points>
<intersection>-71 2</intersection>
<intersection>-66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312,-66.5,322,-66.5</points>
<connection>
<GID>168</GID>
<name>IN_6</name></connection>
<intersection>312 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>307.5,-71,312,-71</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>312 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314,-74,314,-67.5</points>
<intersection>-74 2</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-67.5,322,-67.5</points>
<connection>
<GID>168</GID>
<name>IN_5</name></connection>
<intersection>314 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308,-74,314,-74</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>314 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316,-76.5,316,-68.5</points>
<intersection>-76.5 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>316,-68.5,322,-68.5</points>
<connection>
<GID>168</GID>
<name>IN_4</name></connection>
<intersection>316 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308,-76.5,316,-76.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>316 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>329,-65,332.5,-65</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<connection>
<GID>168</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>316.5,-84.5,321.5,-84.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>321.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>321.5,-88,321.5,-84.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>-84.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>308.5,-87,320,-87</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>320 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>320,-89,320,-87</points>
<intersection>-89 8</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>320,-89,321.5,-89</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>320 7</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319,-90,319,-89.5</points>
<intersection>-90 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319,-90,321.5,-90</points>
<connection>
<GID>221</GID>
<name>IN_2</name></connection>
<intersection>319 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>307,-89.5,319,-89.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>319 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-92,309,-91</points>
<intersection>-92 2</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309,-91,321.5,-91</points>
<connection>
<GID>221</GID>
<name>IN_3</name></connection>
<intersection>309 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>307,-92,309,-92</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,-95,310,-92</points>
<intersection>-95 2</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310,-92,321.5,-92</points>
<connection>
<GID>221</GID>
<name>IN_7</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>307,-95,310,-95</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,-97.5,311.5,-93</points>
<intersection>-97.5 2</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311.5,-93,321.5,-93</points>
<connection>
<GID>221</GID>
<name>IN_6</name></connection>
<intersection>311.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>307,-97.5,311.5,-97.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>311.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313.5,-100.5,313.5,-94</points>
<intersection>-100.5 2</intersection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313.5,-94,321.5,-94</points>
<connection>
<GID>221</GID>
<name>IN_5</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>307.5,-100.5,313.5,-100.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315.5,-103,315.5,-95</points>
<intersection>-103 2</intersection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>315.5,-95,321.5,-95</points>
<connection>
<GID>221</GID>
<name>IN_4</name></connection>
<intersection>315.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>307.5,-103,315.5,-103</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>315.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>328.5,-91.5,332,-91.5</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<connection>
<GID>230</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>314.5,-116,323,-116</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>323 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>323,-120,323,-116</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>-116 1</intersection></vsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>310,-119,321.5,-119</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>321.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>321.5,-121,321.5,-119</points>
<intersection>-121 8</intersection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>321.5,-121,323,-121</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<intersection>321.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320.5,-122,320.5,-121.5</points>
<intersection>-122 1</intersection>
<intersection>-121.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,-122,323,-122</points>
<connection>
<GID>231</GID>
<name>IN_2</name></connection>
<intersection>320.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-121.5,320.5,-121.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>320.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,-124,310.5,-123</points>
<intersection>-124 2</intersection>
<intersection>-123 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310.5,-123,323,-123</points>
<connection>
<GID>231</GID>
<name>IN_3</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-124,310.5,-124</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,-127,311.5,-124</points>
<intersection>-127 2</intersection>
<intersection>-124 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311.5,-124,323,-124</points>
<connection>
<GID>231</GID>
<name>IN_7</name></connection>
<intersection>311.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-127,311.5,-127</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>311.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313,-129.5,313,-125</points>
<intersection>-129.5 2</intersection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313,-125,323,-125</points>
<connection>
<GID>231</GID>
<name>IN_6</name></connection>
<intersection>313 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-129.5,313,-129.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>313 0</intersection></hsegment></shape></wire>
<wire>
<ID>1004</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452,-65.5,452,-61</points>
<intersection>-65.5 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>452,-61,462,-61</points>
<connection>
<GID>991</GID>
<name>IN_6</name></connection>
<intersection>452 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-65.5,452,-65.5</points>
<connection>
<GID>1003</GID>
<name>IN_0</name></connection>
<intersection>452 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315,-132.5,315,-126</points>
<intersection>-132.5 2</intersection>
<intersection>-126 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>315,-126,323,-126</points>
<connection>
<GID>231</GID>
<name>IN_5</name></connection>
<intersection>315 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309,-132.5,315,-132.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>315 0</intersection></hsegment></shape></wire>
<wire>
<ID>1005</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454,-68.5,454,-62</points>
<intersection>-68.5 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>454,-62,462,-62</points>
<connection>
<GID>991</GID>
<name>IN_5</name></connection>
<intersection>454 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448,-68.5,454,-68.5</points>
<connection>
<GID>1004</GID>
<name>IN_0</name></connection>
<intersection>454 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317,-135,317,-127</points>
<intersection>-135 2</intersection>
<intersection>-127 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317,-127,323,-127</points>
<connection>
<GID>231</GID>
<name>IN_4</name></connection>
<intersection>317 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309,-135,317,-135</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>317 0</intersection></hsegment></shape></wire>
<wire>
<ID>1006</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,-71,456,-63</points>
<intersection>-71 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>456,-63,462,-63</points>
<connection>
<GID>991</GID>
<name>IN_4</name></connection>
<intersection>456 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448,-71,456,-71</points>
<connection>
<GID>1005</GID>
<name>IN_0</name></connection>
<intersection>456 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>330,-123.5,333.5,-123.5</points>
<connection>
<GID>231</GID>
<name>OUT</name></connection>
<connection>
<GID>240</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1007</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>469,-59.5,472.5,-59.5</points>
<connection>
<GID>991</GID>
<name>OUT</name></connection>
<connection>
<GID>1006</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>317.5,-139,322.5,-139</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>322.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>322.5,-142.5,322.5,-139</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>-139 1</intersection></vsegment></shape></wire>
<wire>
<ID>1008</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>457,-84,462,-84</points>
<connection>
<GID>1008</GID>
<name>IN_0</name></connection>
<intersection>462 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>462,-87.5,462,-84</points>
<connection>
<GID>1007</GID>
<name>IN_0</name></connection>
<intersection>-84 1</intersection></vsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>309.5,-141.5,321,-141.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>321 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>321,-143.5,321,-141.5</points>
<intersection>-143.5 8</intersection>
<intersection>-141.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>321,-143.5,322.5,-143.5</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>321 7</intersection></hsegment></shape></wire>
<wire>
<ID>1009</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>449,-86.5,460.5,-86.5</points>
<connection>
<GID>1009</GID>
<name>IN_0</name></connection>
<intersection>460.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>460.5,-88.5,460.5,-86.5</points>
<intersection>-88.5 8</intersection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>460.5,-88.5,462,-88.5</points>
<connection>
<GID>1007</GID>
<name>IN_1</name></connection>
<intersection>460.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320,-144.5,320,-144</points>
<intersection>-144.5 1</intersection>
<intersection>-144 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320,-144.5,322.5,-144.5</points>
<connection>
<GID>242</GID>
<name>IN_2</name></connection>
<intersection>320 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308,-144,320,-144</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>320 0</intersection></hsegment></shape></wire>
<wire>
<ID>1010</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459.5,-89.5,459.5,-89</points>
<intersection>-89.5 1</intersection>
<intersection>-89 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>459.5,-89.5,462,-89.5</points>
<connection>
<GID>1007</GID>
<name>IN_2</name></connection>
<intersection>459.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-89,459.5,-89</points>
<connection>
<GID>1010</GID>
<name>IN_0</name></connection>
<intersection>459.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,-146.5,310,-145.5</points>
<intersection>-146.5 2</intersection>
<intersection>-145.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310,-145.5,322.5,-145.5</points>
<connection>
<GID>242</GID>
<name>IN_3</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308,-146.5,310,-146.5</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>1011</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449.5,-91.5,449.5,-90.5</points>
<intersection>-91.5 2</intersection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>449.5,-90.5,462,-90.5</points>
<connection>
<GID>1007</GID>
<name>IN_3</name></connection>
<intersection>449.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-91.5,449.5,-91.5</points>
<connection>
<GID>1011</GID>
<name>IN_0</name></connection>
<intersection>449.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-149.5,311,-146.5</points>
<intersection>-149.5 2</intersection>
<intersection>-146.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311,-146.5,322.5,-146.5</points>
<connection>
<GID>242</GID>
<name>IN_7</name></connection>
<intersection>311 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308,-149.5,311,-149.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>311 0</intersection></hsegment></shape></wire>
<wire>
<ID>1012</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>450.5,-94.5,450.5,-91.5</points>
<intersection>-94.5 2</intersection>
<intersection>-91.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>450.5,-91.5,462,-91.5</points>
<connection>
<GID>1007</GID>
<name>IN_7</name></connection>
<intersection>450.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-94.5,450.5,-94.5</points>
<connection>
<GID>1012</GID>
<name>IN_0</name></connection>
<intersection>450.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312.5,-152,312.5,-147.5</points>
<intersection>-152 2</intersection>
<intersection>-147.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312.5,-147.5,322.5,-147.5</points>
<connection>
<GID>242</GID>
<name>IN_6</name></connection>
<intersection>312.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308,-152,312.5,-152</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>312.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1013</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452,-97,452,-92.5</points>
<intersection>-97 2</intersection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>452,-92.5,462,-92.5</points>
<connection>
<GID>1007</GID>
<name>IN_6</name></connection>
<intersection>452 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-97,452,-97</points>
<connection>
<GID>1013</GID>
<name>IN_0</name></connection>
<intersection>452 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314.5,-155,314.5,-148.5</points>
<intersection>-155 2</intersection>
<intersection>-148.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314.5,-148.5,322.5,-148.5</points>
<connection>
<GID>242</GID>
<name>IN_5</name></connection>
<intersection>314.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-155,314.5,-155</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>314.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1014</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454,-100,454,-93.5</points>
<intersection>-100 2</intersection>
<intersection>-93.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>454,-93.5,462,-93.5</points>
<connection>
<GID>1007</GID>
<name>IN_5</name></connection>
<intersection>454 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448,-100,454,-100</points>
<connection>
<GID>1014</GID>
<name>IN_0</name></connection>
<intersection>454 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316.5,-157.5,316.5,-149.5</points>
<intersection>-157.5 2</intersection>
<intersection>-149.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>316.5,-149.5,322.5,-149.5</points>
<connection>
<GID>242</GID>
<name>IN_4</name></connection>
<intersection>316.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-157.5,316.5,-157.5</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>316.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1015</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,-102.5,456,-94.5</points>
<intersection>-102.5 2</intersection>
<intersection>-94.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>456,-94.5,462,-94.5</points>
<connection>
<GID>1007</GID>
<name>IN_4</name></connection>
<intersection>456 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448,-102.5,456,-102.5</points>
<connection>
<GID>1015</GID>
<name>IN_0</name></connection>
<intersection>456 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>329.5,-146,333,-146</points>
<connection>
<GID>242</GID>
<name>OUT</name></connection>
<connection>
<GID>251</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1016</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>469,-91,472.5,-91</points>
<connection>
<GID>1007</GID>
<name>OUT</name></connection>
<connection>
<GID>1016</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-184,128,-184</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>128 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128,-187.5,128,-184</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>-184 1</intersection></vsegment></shape></wire>
<wire>
<ID>1017</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>460,-150,465,-150</points>
<connection>
<GID>1018</GID>
<name>IN_0</name></connection>
<intersection>465 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>465,-153.5,465,-150</points>
<connection>
<GID>1017</GID>
<name>IN_0</name></connection>
<intersection>-150 1</intersection></vsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115,-186.5,126.5,-186.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>126.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>126.5,-188.5,126.5,-186.5</points>
<intersection>-188.5 8</intersection>
<intersection>-186.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>126.5,-188.5,128,-188.5</points>
<connection>
<GID>252</GID>
<name>IN_1</name></connection>
<intersection>126.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1018</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>452,-152.5,463.5,-152.5</points>
<connection>
<GID>1019</GID>
<name>IN_0</name></connection>
<intersection>463.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>463.5,-154.5,463.5,-152.5</points>
<intersection>-154.5 8</intersection>
<intersection>-152.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>463.5,-154.5,465,-154.5</points>
<connection>
<GID>1017</GID>
<name>IN_1</name></connection>
<intersection>463.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-189.5,125.5,-189</points>
<intersection>-189.5 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125.5,-189.5,128,-189.5</points>
<connection>
<GID>252</GID>
<name>IN_2</name></connection>
<intersection>125.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-189,125.5,-189</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1019</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462.5,-155.5,462.5,-155</points>
<intersection>-155.5 1</intersection>
<intersection>-155 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>462.5,-155.5,465,-155.5</points>
<connection>
<GID>1017</GID>
<name>IN_2</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450.5,-155,462.5,-155</points>
<connection>
<GID>1020</GID>
<name>IN_0</name></connection>
<intersection>462.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-191.5,115.5,-190.5</points>
<intersection>-191.5 2</intersection>
<intersection>-190.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-190.5,128,-190.5</points>
<connection>
<GID>252</GID>
<name>IN_3</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-191.5,115.5,-191.5</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1020</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452.5,-157.5,452.5,-156.5</points>
<intersection>-157.5 2</intersection>
<intersection>-156.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>452.5,-156.5,465,-156.5</points>
<connection>
<GID>1017</GID>
<name>IN_3</name></connection>
<intersection>452.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450.5,-157.5,452.5,-157.5</points>
<connection>
<GID>1021</GID>
<name>IN_0</name></connection>
<intersection>452.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-194.5,116.5,-191.5</points>
<intersection>-194.5 2</intersection>
<intersection>-191.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-191.5,128,-191.5</points>
<connection>
<GID>252</GID>
<name>IN_7</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-194.5,116.5,-194.5</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1021</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>453.5,-160.5,453.5,-157.5</points>
<intersection>-160.5 2</intersection>
<intersection>-157.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>453.5,-157.5,465,-157.5</points>
<connection>
<GID>1017</GID>
<name>IN_7</name></connection>
<intersection>453.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450.5,-160.5,453.5,-160.5</points>
<connection>
<GID>1022</GID>
<name>IN_0</name></connection>
<intersection>453.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-197,118,-192.5</points>
<intersection>-197 2</intersection>
<intersection>-192.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-192.5,128,-192.5</points>
<connection>
<GID>252</GID>
<name>IN_6</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-197,118,-197</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>1022</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455,-163,455,-158.5</points>
<intersection>-163 2</intersection>
<intersection>-158.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>455,-158.5,465,-158.5</points>
<connection>
<GID>1017</GID>
<name>IN_6</name></connection>
<intersection>455 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450.5,-163,455,-163</points>
<connection>
<GID>1023</GID>
<name>IN_0</name></connection>
<intersection>455 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-200,120,-193.5</points>
<intersection>-200 2</intersection>
<intersection>-193.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-193.5,128,-193.5</points>
<connection>
<GID>252</GID>
<name>IN_5</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-200,120,-200</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>1023</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457,-166,457,-159.5</points>
<intersection>-166 2</intersection>
<intersection>-159.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>457,-159.5,465,-159.5</points>
<connection>
<GID>1017</GID>
<name>IN_5</name></connection>
<intersection>457 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>451,-166,457,-166</points>
<connection>
<GID>1024</GID>
<name>IN_0</name></connection>
<intersection>457 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-202.5,122,-194.5</points>
<intersection>-202.5 2</intersection>
<intersection>-194.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,-194.5,128,-194.5</points>
<connection>
<GID>252</GID>
<name>IN_4</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-202.5,122,-202.5</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>1024</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459,-168.5,459,-160.5</points>
<intersection>-168.5 2</intersection>
<intersection>-160.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>459,-160.5,465,-160.5</points>
<connection>
<GID>1017</GID>
<name>IN_4</name></connection>
<intersection>459 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>451,-168.5,459,-168.5</points>
<connection>
<GID>1025</GID>
<name>IN_0</name></connection>
<intersection>459 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135,-191,138.5,-191</points>
<connection>
<GID>252</GID>
<name>OUT</name></connection>
<connection>
<GID>262</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1025</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>472,-157,475.5,-157</points>
<connection>
<GID>1017</GID>
<name>OUT</name></connection>
<connection>
<GID>1026</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1026</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>460,-176,465,-176</points>
<connection>
<GID>1028</GID>
<name>IN_0</name></connection>
<intersection>465 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>465,-179.5,465,-176</points>
<connection>
<GID>1027</GID>
<name>IN_0</name></connection>
<intersection>-176 1</intersection></vsegment></shape></wire>
<wire>
<ID>1027</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>452,-178.5,463.5,-178.5</points>
<connection>
<GID>1029</GID>
<name>IN_0</name></connection>
<intersection>463.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>463.5,-180.5,463.5,-178.5</points>
<intersection>-180.5 8</intersection>
<intersection>-178.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>463.5,-180.5,465,-180.5</points>
<connection>
<GID>1027</GID>
<name>IN_1</name></connection>
<intersection>463.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1028</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462.5,-181.5,462.5,-181</points>
<intersection>-181.5 1</intersection>
<intersection>-181 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>462.5,-181.5,465,-181.5</points>
<connection>
<GID>1027</GID>
<name>IN_2</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450.5,-181,462.5,-181</points>
<connection>
<GID>1030</GID>
<name>IN_0</name></connection>
<intersection>462.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1029</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452.5,-183.5,452.5,-182.5</points>
<intersection>-183.5 2</intersection>
<intersection>-182.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>452.5,-182.5,465,-182.5</points>
<connection>
<GID>1027</GID>
<name>IN_3</name></connection>
<intersection>452.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450.5,-183.5,452.5,-183.5</points>
<connection>
<GID>1031</GID>
<name>IN_0</name></connection>
<intersection>452.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>318,-161,323,-161</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>323 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>323,-164.5,323,-161</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>-161 1</intersection></vsegment></shape></wire>
<wire>
<ID>1030</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>453.5,-186.5,453.5,-183.5</points>
<intersection>-186.5 2</intersection>
<intersection>-183.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>453.5,-183.5,465,-183.5</points>
<connection>
<GID>1027</GID>
<name>IN_7</name></connection>
<intersection>453.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450.5,-186.5,453.5,-186.5</points>
<connection>
<GID>1032</GID>
<name>IN_0</name></connection>
<intersection>453.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>310,-163.5,321.5,-163.5</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>321.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>321.5,-165.5,321.5,-163.5</points>
<intersection>-165.5 8</intersection>
<intersection>-163.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>321.5,-165.5,323,-165.5</points>
<connection>
<GID>280</GID>
<name>IN_1</name></connection>
<intersection>321.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1031</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455,-189,455,-184.5</points>
<intersection>-189 2</intersection>
<intersection>-184.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>455,-184.5,465,-184.5</points>
<connection>
<GID>1027</GID>
<name>IN_6</name></connection>
<intersection>455 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450.5,-189,455,-189</points>
<connection>
<GID>1033</GID>
<name>IN_0</name></connection>
<intersection>455 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320.5,-166.5,320.5,-166</points>
<intersection>-166.5 1</intersection>
<intersection>-166 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,-166.5,323,-166.5</points>
<connection>
<GID>280</GID>
<name>IN_2</name></connection>
<intersection>320.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-166,320.5,-166</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>320.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1032</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457,-192,457,-185.5</points>
<intersection>-192 2</intersection>
<intersection>-185.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>457,-185.5,465,-185.5</points>
<connection>
<GID>1027</GID>
<name>IN_5</name></connection>
<intersection>457 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>451,-192,457,-192</points>
<connection>
<GID>1034</GID>
<name>IN_0</name></connection>
<intersection>457 0</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,-168.5,310.5,-167.5</points>
<intersection>-168.5 2</intersection>
<intersection>-167.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310.5,-167.5,323,-167.5</points>
<connection>
<GID>280</GID>
<name>IN_3</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-168.5,310.5,-168.5</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1033</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459,-194.5,459,-186.5</points>
<intersection>-194.5 2</intersection>
<intersection>-186.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>459,-186.5,465,-186.5</points>
<connection>
<GID>1027</GID>
<name>IN_4</name></connection>
<intersection>459 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>451,-194.5,459,-194.5</points>
<connection>
<GID>1035</GID>
<name>IN_0</name></connection>
<intersection>459 0</intersection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,-171.5,311.5,-168.5</points>
<intersection>-171.5 2</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311.5,-168.5,323,-168.5</points>
<connection>
<GID>280</GID>
<name>IN_7</name></connection>
<intersection>311.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-171.5,311.5,-171.5</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>311.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1034</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>472,-183,475.5,-183</points>
<connection>
<GID>1027</GID>
<name>OUT</name></connection>
<connection>
<GID>1036</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313,-174,313,-169.5</points>
<intersection>-174 2</intersection>
<intersection>-169.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313,-169.5,323,-169.5</points>
<connection>
<GID>280</GID>
<name>IN_6</name></connection>
<intersection>313 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-174,313,-174</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>313 0</intersection></hsegment></shape></wire>
<wire>
<ID>1035</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>457,-206,462,-206</points>
<connection>
<GID>1038</GID>
<name>IN_0</name></connection>
<intersection>462 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>462,-209.5,462,-206</points>
<connection>
<GID>1037</GID>
<name>IN_0</name></connection>
<intersection>-206 1</intersection></vsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315,-177,315,-170.5</points>
<intersection>-177 2</intersection>
<intersection>-170.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>315,-170.5,323,-170.5</points>
<connection>
<GID>280</GID>
<name>IN_5</name></connection>
<intersection>315 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309,-177,315,-177</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>315 0</intersection></hsegment></shape></wire>
<wire>
<ID>1036</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>449,-208.5,460.5,-208.5</points>
<connection>
<GID>1039</GID>
<name>IN_0</name></connection>
<intersection>460.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>460.5,-210.5,460.5,-208.5</points>
<intersection>-210.5 8</intersection>
<intersection>-208.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>460.5,-210.5,462,-210.5</points>
<connection>
<GID>1037</GID>
<name>IN_1</name></connection>
<intersection>460.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317,-179.5,317,-171.5</points>
<intersection>-179.5 2</intersection>
<intersection>-171.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317,-171.5,323,-171.5</points>
<connection>
<GID>280</GID>
<name>IN_4</name></connection>
<intersection>317 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309,-179.5,317,-179.5</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>317 0</intersection></hsegment></shape></wire>
<wire>
<ID>1037</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459.5,-211.5,459.5,-211</points>
<intersection>-211.5 1</intersection>
<intersection>-211 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>459.5,-211.5,462,-211.5</points>
<connection>
<GID>1037</GID>
<name>IN_2</name></connection>
<intersection>459.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-211,459.5,-211</points>
<connection>
<GID>1040</GID>
<name>IN_0</name></connection>
<intersection>459.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>330,-168,333.5,-168</points>
<connection>
<GID>280</GID>
<name>OUT</name></connection>
<connection>
<GID>289</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1038</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449.5,-213.5,449.5,-212.5</points>
<intersection>-213.5 2</intersection>
<intersection>-212.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>449.5,-212.5,462,-212.5</points>
<connection>
<GID>1037</GID>
<name>IN_3</name></connection>
<intersection>449.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-213.5,449.5,-213.5</points>
<connection>
<GID>1041</GID>
<name>IN_0</name></connection>
<intersection>449.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1039</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>450.5,-216.5,450.5,-213.5</points>
<intersection>-216.5 2</intersection>
<intersection>-213.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>450.5,-213.5,462,-213.5</points>
<connection>
<GID>1037</GID>
<name>IN_7</name></connection>
<intersection>450.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-216.5,450.5,-216.5</points>
<connection>
<GID>1042</GID>
<name>IN_0</name></connection>
<intersection>450.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1040</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452,-219,452,-214.5</points>
<intersection>-219 2</intersection>
<intersection>-214.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>452,-214.5,462,-214.5</points>
<connection>
<GID>1037</GID>
<name>IN_6</name></connection>
<intersection>452 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-219,452,-219</points>
<connection>
<GID>1043</GID>
<name>IN_0</name></connection>
<intersection>452 0</intersection></hsegment></shape></wire>
<wire>
<ID>1041</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>454,-222,454,-215.5</points>
<intersection>-222 2</intersection>
<intersection>-215.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>454,-215.5,462,-215.5</points>
<connection>
<GID>1037</GID>
<name>IN_5</name></connection>
<intersection>454 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448,-222,454,-222</points>
<connection>
<GID>1044</GID>
<name>IN_0</name></connection>
<intersection>454 0</intersection></hsegment></shape></wire>
<wire>
<ID>1042</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,-224.5,456,-216.5</points>
<intersection>-224.5 2</intersection>
<intersection>-216.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>456,-216.5,462,-216.5</points>
<connection>
<GID>1037</GID>
<name>IN_4</name></connection>
<intersection>456 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448,-224.5,456,-224.5</points>
<connection>
<GID>1045</GID>
<name>IN_0</name></connection>
<intersection>456 0</intersection></hsegment></shape></wire>
<wire>
<ID>1043</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>469,-213,472.5,-213</points>
<connection>
<GID>1037</GID>
<name>OUT</name></connection>
<connection>
<GID>1046</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1044</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>456.5,-230.5,461.5,-230.5</points>
<connection>
<GID>1048</GID>
<name>IN_0</name></connection>
<intersection>461.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>461.5,-234,461.5,-230.5</points>
<connection>
<GID>1047</GID>
<name>IN_0</name></connection>
<intersection>-230.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1045</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>448.5,-233,460,-233</points>
<connection>
<GID>1049</GID>
<name>IN_0</name></connection>
<intersection>460 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>460,-235,460,-233</points>
<intersection>-235 8</intersection>
<intersection>-233 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>460,-235,461.5,-235</points>
<connection>
<GID>1047</GID>
<name>IN_1</name></connection>
<intersection>460 7</intersection></hsegment></shape></wire>
<wire>
<ID>1046</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459,-236,459,-235.5</points>
<intersection>-236 1</intersection>
<intersection>-235.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>459,-236,461.5,-236</points>
<connection>
<GID>1047</GID>
<name>IN_2</name></connection>
<intersection>459 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447,-235.5,459,-235.5</points>
<connection>
<GID>1050</GID>
<name>IN_0</name></connection>
<intersection>459 0</intersection></hsegment></shape></wire>
<wire>
<ID>1047</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449,-238,449,-237</points>
<intersection>-238 2</intersection>
<intersection>-237 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>449,-237,461.5,-237</points>
<connection>
<GID>1047</GID>
<name>IN_3</name></connection>
<intersection>449 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447,-238,449,-238</points>
<connection>
<GID>1051</GID>
<name>IN_0</name></connection>
<intersection>449 0</intersection></hsegment></shape></wire>
<wire>
<ID>1048</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>450,-241,450,-238</points>
<intersection>-241 2</intersection>
<intersection>-238 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>450,-238,461.5,-238</points>
<connection>
<GID>1047</GID>
<name>IN_7</name></connection>
<intersection>450 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447,-241,450,-241</points>
<connection>
<GID>1052</GID>
<name>IN_0</name></connection>
<intersection>450 0</intersection></hsegment></shape></wire>
<wire>
<ID>1049</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>451.5,-243.5,451.5,-239</points>
<intersection>-243.5 2</intersection>
<intersection>-239 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>451.5,-239,461.5,-239</points>
<connection>
<GID>1047</GID>
<name>IN_6</name></connection>
<intersection>451.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447,-243.5,451.5,-243.5</points>
<connection>
<GID>1053</GID>
<name>IN_0</name></connection>
<intersection>451.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1050</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>453.5,-246.5,453.5,-240</points>
<intersection>-246.5 2</intersection>
<intersection>-240 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>453.5,-240,461.5,-240</points>
<connection>
<GID>1047</GID>
<name>IN_5</name></connection>
<intersection>453.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-246.5,453.5,-246.5</points>
<connection>
<GID>1054</GID>
<name>IN_0</name></connection>
<intersection>453.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1051</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455.5,-249,455.5,-241</points>
<intersection>-249 2</intersection>
<intersection>-241 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>455.5,-241,461.5,-241</points>
<connection>
<GID>1047</GID>
<name>IN_4</name></connection>
<intersection>455.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>447.5,-249,455.5,-249</points>
<connection>
<GID>1055</GID>
<name>IN_0</name></connection>
<intersection>455.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1052</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>468.5,-237.5,472,-237.5</points>
<connection>
<GID>1047</GID>
<name>OUT</name></connection>
<connection>
<GID>1056</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1053</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>509,-52.5,514,-52.5</points>
<connection>
<GID>1060</GID>
<name>IN_0</name></connection>
<intersection>514 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>514,-56,514,-52.5</points>
<connection>
<GID>1059</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1054</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>501,-55,512.5,-55</points>
<connection>
<GID>1061</GID>
<name>IN_0</name></connection>
<intersection>512.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>512.5,-57,512.5,-55</points>
<intersection>-57 8</intersection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>512.5,-57,514,-57</points>
<connection>
<GID>1059</GID>
<name>IN_1</name></connection>
<intersection>512.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1055</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511.5,-58,511.5,-57.5</points>
<intersection>-58 1</intersection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511.5,-58,514,-58</points>
<connection>
<GID>1059</GID>
<name>IN_2</name></connection>
<intersection>511.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>499.5,-57.5,511.5,-57.5</points>
<connection>
<GID>1062</GID>
<name>IN_0</name></connection>
<intersection>511.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1056</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>501.5,-60,501.5,-59</points>
<intersection>-60 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>501.5,-59,514,-59</points>
<connection>
<GID>1059</GID>
<name>IN_3</name></connection>
<intersection>501.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>499.5,-60,501.5,-60</points>
<connection>
<GID>1063</GID>
<name>IN_0</name></connection>
<intersection>501.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1057</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502.5,-63,502.5,-60</points>
<intersection>-63 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>502.5,-60,514,-60</points>
<connection>
<GID>1059</GID>
<name>IN_7</name></connection>
<intersection>502.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>499.5,-63,502.5,-63</points>
<connection>
<GID>1064</GID>
<name>IN_0</name></connection>
<intersection>502.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1058</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>504,-65.5,504,-61</points>
<intersection>-65.5 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>504,-61,514,-61</points>
<connection>
<GID>1059</GID>
<name>IN_6</name></connection>
<intersection>504 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>499.5,-65.5,504,-65.5</points>
<connection>
<GID>1065</GID>
<name>IN_0</name></connection>
<intersection>504 0</intersection></hsegment></shape></wire>
<wire>
<ID>1059</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>506,-68.5,506,-62</points>
<intersection>-68.5 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>506,-62,514,-62</points>
<connection>
<GID>1059</GID>
<name>IN_5</name></connection>
<intersection>506 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>500,-68.5,506,-68.5</points>
<connection>
<GID>1066</GID>
<name>IN_0</name></connection>
<intersection>506 0</intersection></hsegment></shape></wire>
<wire>
<ID>1060</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>508,-71,508,-63</points>
<intersection>-71 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>508,-63,514,-63</points>
<connection>
<GID>1059</GID>
<name>IN_4</name></connection>
<intersection>508 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>500,-71,508,-71</points>
<connection>
<GID>1067</GID>
<name>IN_0</name></connection>
<intersection>508 0</intersection></hsegment></shape></wire>
<wire>
<ID>1061</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>521,-59.5,524.5,-59.5</points>
<connection>
<GID>1059</GID>
<name>OUT</name></connection>
<connection>
<GID>1068</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>705</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-83,170,-83</points>
<connection>
<GID>580</GID>
<name>IN_0</name></connection>
<intersection>170 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>170,-86.5,170,-83</points>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<intersection>-83 1</intersection></vsegment></shape></wire>
<wire>
<ID>706</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-85.5,168.5,-85.5</points>
<connection>
<GID>581</GID>
<name>IN_0</name></connection>
<intersection>168.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>168.5,-87.5,168.5,-85.5</points>
<intersection>-87.5 8</intersection>
<intersection>-85.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>168.5,-87.5,170,-87.5</points>
<connection>
<GID>579</GID>
<name>IN_1</name></connection>
<intersection>168.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>707</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-88.5,167.5,-88</points>
<intersection>-88.5 1</intersection>
<intersection>-88 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167.5,-88.5,170,-88.5</points>
<connection>
<GID>579</GID>
<name>IN_2</name></connection>
<intersection>167.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155.5,-88,167.5,-88</points>
<connection>
<GID>582</GID>
<name>IN_0</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>708</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,-90.5,157.5,-89.5</points>
<intersection>-90.5 2</intersection>
<intersection>-89.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-89.5,170,-89.5</points>
<connection>
<GID>579</GID>
<name>IN_3</name></connection>
<intersection>157.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155.5,-90.5,157.5,-90.5</points>
<connection>
<GID>583</GID>
<name>IN_0</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>709</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158.5,-93.5,158.5,-90.5</points>
<intersection>-93.5 2</intersection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158.5,-90.5,170,-90.5</points>
<connection>
<GID>579</GID>
<name>IN_7</name></connection>
<intersection>158.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155.5,-93.5,158.5,-93.5</points>
<connection>
<GID>584</GID>
<name>IN_0</name></connection>
<intersection>158.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>710</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-96,160,-91.5</points>
<intersection>-96 2</intersection>
<intersection>-91.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160,-91.5,170,-91.5</points>
<connection>
<GID>579</GID>
<name>IN_6</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155.5,-96,160,-96</points>
<connection>
<GID>585</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>711</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-99,162,-92.5</points>
<intersection>-99 2</intersection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162,-92.5,170,-92.5</points>
<connection>
<GID>579</GID>
<name>IN_5</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156,-99,162,-99</points>
<connection>
<GID>587</GID>
<name>IN_0</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>712</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164,-101.5,164,-93.5</points>
<intersection>-101.5 2</intersection>
<intersection>-93.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164,-93.5,170,-93.5</points>
<connection>
<GID>579</GID>
<name>IN_4</name></connection>
<intersection>164 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156,-101.5,164,-101.5</points>
<connection>
<GID>595</GID>
<name>IN_0</name></connection>
<intersection>164 0</intersection></hsegment></shape></wire>
<wire>
<ID>713</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-90,180.5,-90</points>
<connection>
<GID>579</GID>
<name>OUT</name></connection>
<connection>
<GID>598</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,-60,175,-59.5</points>
<intersection>-60 1</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-60,177.5,-60</points>
<connection>
<GID>325</GID>
<name>IN_2</name></connection>
<intersection>175 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163,-59.5,175,-59.5</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>175 0</intersection></hsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-62,165,-61</points>
<intersection>-62 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165,-61,177.5,-61</points>
<connection>
<GID>325</GID>
<name>IN_3</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163,-62,165,-62</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>730</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>319,-191,324,-191</points>
<connection>
<GID>728</GID>
<name>IN_0</name></connection>
<intersection>324 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>324,-194.5,324,-191</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>-191 1</intersection></vsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-65,166,-62</points>
<intersection>-65 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-62,177.5,-62</points>
<connection>
<GID>325</GID>
<name>IN_7</name></connection>
<intersection>166 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163,-65,166,-65</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>731</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>311,-193.5,322.5,-193.5</points>
<connection>
<GID>730</GID>
<name>IN_0</name></connection>
<intersection>322.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>322.5,-195.5,322.5,-193.5</points>
<intersection>-195.5 8</intersection>
<intersection>-193.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>322.5,-195.5,324,-195.5</points>
<connection>
<GID>726</GID>
<name>IN_1</name></connection>
<intersection>322.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-67.5,167.5,-63</points>
<intersection>-67.5 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167.5,-63,177.5,-63</points>
<connection>
<GID>325</GID>
<name>IN_6</name></connection>
<intersection>167.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163,-67.5,167.5,-67.5</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>732</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321.5,-196.5,321.5,-196</points>
<intersection>-196.5 1</intersection>
<intersection>-196 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321.5,-196.5,324,-196.5</points>
<connection>
<GID>726</GID>
<name>IN_2</name></connection>
<intersection>321.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309.5,-196,321.5,-196</points>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<intersection>321.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>733</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,-198.5,311.5,-197.5</points>
<intersection>-198.5 2</intersection>
<intersection>-197.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311.5,-197.5,324,-197.5</points>
<connection>
<GID>726</GID>
<name>IN_3</name></connection>
<intersection>311.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309.5,-198.5,311.5,-198.5</points>
<connection>
<GID>732</GID>
<name>IN_0</name></connection>
<intersection>311.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>734</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312.5,-201.5,312.5,-198.5</points>
<intersection>-201.5 2</intersection>
<intersection>-198.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312.5,-198.5,324,-198.5</points>
<connection>
<GID>726</GID>
<name>IN_7</name></connection>
<intersection>312.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309.5,-201.5,312.5,-201.5</points>
<connection>
<GID>733</GID>
<name>IN_0</name></connection>
<intersection>312.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314,-204,314,-199.5</points>
<intersection>-204 2</intersection>
<intersection>-199.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-199.5,324,-199.5</points>
<connection>
<GID>726</GID>
<name>IN_6</name></connection>
<intersection>314 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309.5,-204,314,-204</points>
<connection>
<GID>738</GID>
<name>IN_0</name></connection>
<intersection>314 0</intersection></hsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316,-207,316,-200.5</points>
<intersection>-207 2</intersection>
<intersection>-200.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>316,-200.5,324,-200.5</points>
<connection>
<GID>726</GID>
<name>IN_5</name></connection>
<intersection>316 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>310,-207,316,-207</points>
<connection>
<GID>742</GID>
<name>IN_0</name></connection>
<intersection>316 0</intersection></hsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318,-209.5,318,-201.5</points>
<intersection>-209.5 2</intersection>
<intersection>-201.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318,-201.5,324,-201.5</points>
<connection>
<GID>726</GID>
<name>IN_4</name></connection>
<intersection>318 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>310,-209.5,318,-209.5</points>
<connection>
<GID>743</GID>
<name>IN_0</name></connection>
<intersection>318 0</intersection></hsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>331,-198,334.5,-198</points>
<connection>
<GID>744</GID>
<name>IN_0</name></connection>
<connection>
<GID>726</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-70.5,169.5,-64</points>
<intersection>-70.5 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-64,177.5,-64</points>
<connection>
<GID>325</GID>
<name>IN_5</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163.5,-70.5,169.5,-70.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171.5,-73,171.5,-65</points>
<intersection>-73 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171.5,-65,177.5,-65</points>
<connection>
<GID>325</GID>
<name>IN_4</name></connection>
<intersection>171.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163.5,-73,171.5,-73</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>171.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>184.5,-61.5,188,-61.5</points>
<connection>
<GID>325</GID>
<name>OUT</name></connection>
<connection>
<GID>334</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-49,163.5,-47.5</points>
<intersection>-49 1</intersection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163.5,-49,165.5,-49</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-47.5,163.5,-47.5</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-51.5,163.5,-51</points>
<intersection>-51.5 2</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163.5,-51,165.5,-51</points>
<connection>
<GID>365</GID>
<name>IN_1</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155.5,-51.5,163.5,-51.5</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<intersection>158 3</intersection>
<intersection>163.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>158,-55,158,-51.5</points>
<intersection>-55 4</intersection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>158,-55,158.5,-55</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>158 3</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-58,174,-50</points>
<intersection>-58 1</intersection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,-58,177.5,-58</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>171.5,-50,174,-50</points>
<connection>
<GID>365</GID>
<name>OUT</name></connection>
<intersection>174 0</intersection></hsegment></shape></wire>
<wire>
<ID>763</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>459.5,-118.5,464.5,-118.5</points>
<connection>
<GID>947</GID>
<name>IN_0</name></connection>
<intersection>464.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>464.5,-122,464.5,-118.5</points>
<connection>
<GID>900</GID>
<name>IN_0</name></connection>
<intersection>-118.5 1</intersection></vsegment></shape></wire></page 3>
<page 4>
<PageViewport>163.693,0.0220676,676.031,-293.913</PageViewport>
<gate>
<ID>389</ID>
<type>GA_LED</type>
<position>-56.5,-4.5</position>
<input>
<ID>N_in2</ID>315 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>390</ID>
<type>DE_TO</type>
<position>-65,-96.5</position>
<input>
<ID>IN_0</ID>661 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A12</lparam></gate>
<gate>
<ID>391</ID>
<type>DE_TO</type>
<position>-70.5,-95</position>
<input>
<ID>IN_0</ID>334 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A13</lparam></gate>
<gate>
<ID>392</ID>
<type>DE_TO</type>
<position>-64,-93.5</position>
<input>
<ID>IN_0</ID>335 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A14</lparam></gate>
<gate>
<ID>393</ID>
<type>DE_TO</type>
<position>-70,-92</position>
<input>
<ID>IN_0</ID>336 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A15</lparam></gate>
<gate>
<ID>394</ID>
<type>DE_TO</type>
<position>-60,-7.5</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Zero</lparam></gate>
<gate>
<ID>395</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>3,-43</position>
<input>
<ID>ENABLE_0</ID>396 </input>
<input>
<ID>IN_0</ID>350 </input>
<input>
<ID>IN_1</ID>349 </input>
<input>
<ID>IN_2</ID>348 </input>
<input>
<ID>IN_3</ID>347 </input>
<output>
<ID>OUT_0</ID>346 </output>
<output>
<ID>OUT_1</ID>345 </output>
<output>
<ID>OUT_2</ID>344 </output>
<output>
<ID>OUT_3</ID>343 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>396</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>6.5,-33.5</position>
<input>
<ID>ENABLE_0</ID>369 </input>
<input>
<ID>IN_0</ID>354 </input>
<input>
<ID>IN_1</ID>353 </input>
<input>
<ID>IN_2</ID>352 </input>
<input>
<ID>IN_3</ID>351 </input>
<output>
<ID>OUT_0</ID>343 </output>
<output>
<ID>OUT_1</ID>344 </output>
<output>
<ID>OUT_2</ID>345 </output>
<output>
<ID>OUT_3</ID>346 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>397</ID>
<type>BE_NOR4</type>
<position>-31.5,-83.5</position>
<input>
<ID>IN_0</ID>661 </input>
<input>
<ID>IN_1</ID>334 </input>
<input>
<ID>IN_2</ID>335 </input>
<input>
<ID>IN_3</ID>336 </input>
<output>
<ID>OUT</ID>418 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>398</ID>
<type>DA_FROM</type>
<position>-4,-41.5</position>
<input>
<ID>IN_0</ID>347 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A15</lparam></gate>
<gate>
<ID>399</ID>
<type>DA_FROM</type>
<position>-8.5,-42.5</position>
<input>
<ID>IN_0</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A14</lparam></gate>
<gate>
<ID>400</ID>
<type>DA_FROM</type>
<position>-14,-43.5</position>
<input>
<ID>IN_0</ID>349 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A13</lparam></gate>
<gate>
<ID>401</ID>
<type>DA_FROM</type>
<position>-20,-44.5</position>
<input>
<ID>IN_0</ID>350 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A12</lparam></gate>
<gate>
<ID>402</ID>
<type>DA_FROM</type>
<position>55,-22.5</position>
<input>
<ID>IN_0</ID>351 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>403</ID>
<type>DA_FROM</type>
<position>51,-22</position>
<input>
<ID>IN_0</ID>352 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>404</ID>
<type>DA_FROM</type>
<position>47,-21.5</position>
<input>
<ID>IN_0</ID>353 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>405</ID>
<type>DA_FROM</type>
<position>44,-21.5</position>
<input>
<ID>IN_0</ID>354 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>406</ID>
<type>DA_FROM</type>
<position>7.5,-49</position>
<input>
<ID>IN_0</ID>355 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>407</ID>
<type>FF_GND</type>
<position>15,-48.5</position>
<output>
<ID>OUT_0</ID>356 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>408</ID>
<type>FF_GND</type>
<position>14,-35.5</position>
<output>
<ID>OUT_0</ID>357 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>409</ID>
<type>DA_FROM</type>
<position>93.5,-22.5</position>
<input>
<ID>IN_0</ID>397 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Res-Acc</lparam></gate>
<gate>
<ID>410</ID>
<type>DA_FROM</type>
<position>183,-29</position>
<input>
<ID>IN_0</ID>398 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Res-Acc</lparam></gate>
<gate>
<ID>411</ID>
<type>DA_FROM</type>
<position>271,-27</position>
<input>
<ID>IN_0</ID>450 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Res-Acc</lparam></gate>
<gate>
<ID>418</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>93.5,-42</position>
<input>
<ID>ENABLE_0</ID>397 </input>
<input>
<ID>IN_0</ID>406 </input>
<input>
<ID>IN_1</ID>405 </input>
<input>
<ID>IN_2</ID>404 </input>
<input>
<ID>IN_3</ID>403 </input>
<output>
<ID>OUT_0</ID>402 </output>
<output>
<ID>OUT_1</ID>401 </output>
<output>
<ID>OUT_2</ID>400 </output>
<output>
<ID>OUT_3</ID>399 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>419</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>97,-32.5</position>
<input>
<ID>ENABLE_0</ID>370 </input>
<input>
<ID>IN_0</ID>410 </input>
<input>
<ID>IN_1</ID>409 </input>
<input>
<ID>IN_2</ID>408 </input>
<input>
<ID>IN_3</ID>407 </input>
<output>
<ID>OUT_0</ID>399 </output>
<output>
<ID>OUT_1</ID>400 </output>
<output>
<ID>OUT_2</ID>401 </output>
<output>
<ID>OUT_3</ID>402 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>420</ID>
<type>DA_FROM</type>
<position>86.5,-40.5</position>
<input>
<ID>IN_0</ID>403 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A11</lparam></gate>
<gate>
<ID>421</ID>
<type>DA_FROM</type>
<position>82,-41.5</position>
<input>
<ID>IN_0</ID>404 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A10</lparam></gate>
<gate>
<ID>422</ID>
<type>DA_FROM</type>
<position>76.5,-42.5</position>
<input>
<ID>IN_0</ID>405 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A9</lparam></gate>
<gate>
<ID>423</ID>
<type>DA_FROM</type>
<position>70.5,-43.5</position>
<input>
<ID>IN_0</ID>406 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A8</lparam></gate>
<gate>
<ID>424</ID>
<type>DA_FROM</type>
<position>148,-22.5</position>
<input>
<ID>IN_0</ID>407 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>425</ID>
<type>DA_FROM</type>
<position>144,-22</position>
<input>
<ID>IN_0</ID>408 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>426</ID>
<type>DA_FROM</type>
<position>140,-21.5</position>
<input>
<ID>IN_0</ID>409 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>427</ID>
<type>DA_FROM</type>
<position>137,-21.5</position>
<input>
<ID>IN_0</ID>410 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>428</ID>
<type>DA_FROM</type>
<position>98,-48</position>
<input>
<ID>IN_0</ID>411 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>429</ID>
<type>FF_GND</type>
<position>105.5,-47.5</position>
<output>
<ID>OUT_0</ID>412 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>430</ID>
<type>FF_GND</type>
<position>104.5,-35</position>
<output>
<ID>OUT_0</ID>413 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>431</ID>
<type>AE_FULLADDER_4BIT</type>
<position>110,-87</position>
<input>
<ID>IN_0</ID>380 </input>
<input>
<ID>IN_1</ID>382 </input>
<input>
<ID>IN_2</ID>383 </input>
<input>
<ID>IN_3</ID>384 </input>
<input>
<ID>IN_B_0</ID>362 </input>
<input>
<ID>IN_B_1</ID>363 </input>
<input>
<ID>IN_B_2</ID>364 </input>
<input>
<ID>IN_B_3</ID>365 </input>
<output>
<ID>OUT_0</ID>390 </output>
<output>
<ID>OUT_1</ID>391 </output>
<output>
<ID>OUT_2</ID>392 </output>
<output>
<ID>OUT_3</ID>393 </output>
<input>
<ID>carry_in</ID>523 </input>
<output>
<ID>carry_out</ID>414 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>432</ID>
<type>AI_XOR2</type>
<position>131,-65.5</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>375 </input>
<output>
<ID>OUT</ID>362 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>433</ID>
<type>AI_XOR2</type>
<position>124.5,-65.5</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>376 </input>
<output>
<ID>OUT</ID>363 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>434</ID>
<type>AI_XOR2</type>
<position>119,-65.5</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>377 </input>
<output>
<ID>OUT</ID>364 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>435</ID>
<type>AI_XOR2</type>
<position>112,-65.5</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>378 </input>
<output>
<ID>OUT</ID>365 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>436</ID>
<type>DA_FROM</type>
<position>106,-58.5</position>
<input>
<ID>IN_0</ID>374 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>437</ID>
<type>DA_FROM</type>
<position>99.5,-58</position>
<input>
<ID>IN_0</ID>373 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>438</ID>
<type>DA_FROM</type>
<position>94.5,-57.5</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>439</ID>
<type>DA_FROM</type>
<position>88,-57.5</position>
<input>
<ID>IN_0</ID>371 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>440</ID>
<type>AI_XOR2</type>
<position>107,-66.5</position>
<input>
<ID>IN_0</ID>388 </input>
<input>
<ID>IN_1</ID>374 </input>
<output>
<ID>OUT</ID>379 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>441</ID>
<type>AI_XOR2</type>
<position>100.5,-66.5</position>
<input>
<ID>IN_0</ID>388 </input>
<input>
<ID>IN_1</ID>373 </input>
<output>
<ID>OUT</ID>381 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>442</ID>
<type>AI_XOR2</type>
<position>95.5,-66.5</position>
<input>
<ID>IN_0</ID>388 </input>
<input>
<ID>IN_1</ID>372 </input>
<output>
<ID>OUT</ID>385 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>443</ID>
<type>AI_XOR2</type>
<position>89,-66.5</position>
<input>
<ID>IN_0</ID>388 </input>
<input>
<ID>IN_1</ID>371 </input>
<output>
<ID>OUT</ID>386 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>450</ID>
<type>AA_REGISTER4</type>
<position>104.5,-42.5</position>
<input>
<ID>IN_0</ID>402 </input>
<input>
<ID>IN_1</ID>401 </input>
<input>
<ID>IN_2</ID>400 </input>
<input>
<ID>IN_3</ID>399 </input>
<output>
<ID>OUT_0</ID>375 </output>
<output>
<ID>OUT_1</ID>376 </output>
<output>
<ID>OUT_2</ID>377 </output>
<output>
<ID>OUT_3</ID>378 </output>
<input>
<ID>clear</ID>412 </input>
<input>
<ID>clock</ID>411 </input>
<input>
<ID>count_enable</ID>413 </input>
<input>
<ID>count_up</ID>413 </input>
<input>
<ID>load</ID>415 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>451</ID>
<type>AA_AND2</type>
<position>108,-75</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>380 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>452</ID>
<type>AA_AND2</type>
<position>101.5,-75.5</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>381 </input>
<output>
<ID>OUT</ID>382 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>453</ID>
<type>AA_AND2</type>
<position>96.5,-75.5</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>385 </input>
<output>
<ID>OUT</ID>383 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>454</ID>
<type>AA_AND2</type>
<position>90,-75.5</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>386 </input>
<output>
<ID>OUT</ID>384 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>455</ID>
<type>AE_SMALL_INVERTER</type>
<position>85.5,-71</position>
<input>
<ID>IN_0</ID>416 </input>
<output>
<ID>OUT_0</ID>387 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>462</ID>
<type>DA_FROM</type>
<position>114.5,-33.5</position>
<input>
<ID>IN_0</ID>415 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LD Acc</lparam></gate>
<gate>
<ID>464</ID>
<type>DA_FROM</type>
<position>76.5,-71</position>
<input>
<ID>IN_0</ID>416 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZero</lparam></gate>
<gate>
<ID>465</ID>
<type>DA_FROM</type>
<position>-11.5,-68.5</position>
<input>
<ID>IN_0</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZero</lparam></gate>
<gate>
<ID>467</ID>
<type>DE_TO</type>
<position>-31.5,-61</position>
<input>
<ID>IN_0</ID>418 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z15-12</lparam></gate>
<gate>
<ID>471</ID>
<type>DA_FROM</type>
<position>-59.5,-36</position>
<input>
<ID>IN_0</ID>624 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z15-12</lparam></gate>
<gate>
<ID>472</ID>
<type>DA_FROM</type>
<position>-56.5,-36</position>
<input>
<ID>IN_0</ID>625 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z11-8</lparam></gate>
<gate>
<ID>475</ID>
<type>DE_TO</type>
<position>58.5,-95.5</position>
<input>
<ID>IN_0</ID>390 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A8</lparam></gate>
<gate>
<ID>476</ID>
<type>DE_TO</type>
<position>53,-94</position>
<input>
<ID>IN_0</ID>391 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A9</lparam></gate>
<gate>
<ID>477</ID>
<type>DE_TO</type>
<position>59.5,-92.5</position>
<input>
<ID>IN_0</ID>392 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A10</lparam></gate>
<gate>
<ID>478</ID>
<type>DE_TO</type>
<position>53.5,-91</position>
<input>
<ID>IN_0</ID>393 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A11</lparam></gate>
<gate>
<ID>479</ID>
<type>DE_TO</type>
<position>287,0</position>
<input>
<ID>IN_0</ID>719 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Ck1</lparam></gate>
<gate>
<ID>480</ID>
<type>BE_NOR4</type>
<position>65.5,-82</position>
<input>
<ID>IN_0</ID>393 </input>
<input>
<ID>IN_1</ID>392 </input>
<input>
<ID>IN_2</ID>391 </input>
<input>
<ID>IN_3</ID>390 </input>
<output>
<ID>OUT</ID>422 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>482</ID>
<type>DE_TO</type>
<position>65.5,-71</position>
<input>
<ID>IN_0</ID>422 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z11-8</lparam></gate>
<gate>
<ID>485</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>183,-42</position>
<input>
<ID>ENABLE_0</ID>398 </input>
<input>
<ID>IN_0</ID>462 </input>
<input>
<ID>IN_1</ID>461 </input>
<input>
<ID>IN_2</ID>460 </input>
<input>
<ID>IN_3</ID>459 </input>
<output>
<ID>OUT_0</ID>458 </output>
<output>
<ID>OUT_1</ID>457 </output>
<output>
<ID>OUT_2</ID>456 </output>
<output>
<ID>OUT_3</ID>455 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>486</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>186.5,-32.5</position>
<input>
<ID>ENABLE_0</ID>394 </input>
<input>
<ID>IN_0</ID>466 </input>
<input>
<ID>IN_1</ID>465 </input>
<input>
<ID>IN_2</ID>464 </input>
<input>
<ID>IN_3</ID>463 </input>
<output>
<ID>OUT_0</ID>455 </output>
<output>
<ID>OUT_1</ID>456 </output>
<output>
<ID>OUT_2</ID>457 </output>
<output>
<ID>OUT_3</ID>458 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>487</ID>
<type>DA_FROM</type>
<position>176,-40.5</position>
<input>
<ID>IN_0</ID>459 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A7</lparam></gate>
<gate>
<ID>488</ID>
<type>DA_FROM</type>
<position>171.5,-41.5</position>
<input>
<ID>IN_0</ID>460 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A6</lparam></gate>
<gate>
<ID>489</ID>
<type>DA_FROM</type>
<position>166,-42.5</position>
<input>
<ID>IN_0</ID>461 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A5</lparam></gate>
<gate>
<ID>490</ID>
<type>DA_FROM</type>
<position>160,-43.5</position>
<input>
<ID>IN_0</ID>462 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A4</lparam></gate>
<gate>
<ID>491</ID>
<type>DA_FROM</type>
<position>235.5,-24.5</position>
<input>
<ID>IN_0</ID>463 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>492</ID>
<type>DA_FROM</type>
<position>231.5,-24</position>
<input>
<ID>IN_0</ID>464 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>493</ID>
<type>DA_FROM</type>
<position>227.5,-23.5</position>
<input>
<ID>IN_0</ID>465 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>494</ID>
<type>DA_FROM</type>
<position>224.5,-23.5</position>
<input>
<ID>IN_0</ID>466 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>495</ID>
<type>DA_FROM</type>
<position>187.5,-48</position>
<input>
<ID>IN_0</ID>467 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>496</ID>
<type>FF_GND</type>
<position>195,-47.5</position>
<output>
<ID>OUT_0</ID>468 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>497</ID>
<type>FF_GND</type>
<position>194,-36</position>
<output>
<ID>OUT_0</ID>469 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>498</ID>
<type>AE_FULLADDER_4BIT</type>
<position>199.5,-87</position>
<input>
<ID>IN_0</ID>436 </input>
<input>
<ID>IN_1</ID>438 </input>
<input>
<ID>IN_2</ID>439 </input>
<input>
<ID>IN_3</ID>440 </input>
<input>
<ID>IN_B_0</ID>423 </input>
<input>
<ID>IN_B_1</ID>424 </input>
<input>
<ID>IN_B_2</ID>425 </input>
<input>
<ID>IN_B_3</ID>426 </input>
<output>
<ID>OUT_0</ID>446 </output>
<output>
<ID>OUT_1</ID>447 </output>
<output>
<ID>OUT_2</ID>448 </output>
<output>
<ID>OUT_3</ID>449 </output>
<input>
<ID>carry_in</ID>524 </input>
<output>
<ID>carry_out</ID>523 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>499</ID>
<type>AI_XOR2</type>
<position>220.5,-65.5</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>431 </input>
<output>
<ID>OUT</ID>423 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>500</ID>
<type>AI_XOR2</type>
<position>214,-65.5</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>432 </input>
<output>
<ID>OUT</ID>424 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>501</ID>
<type>AI_XOR2</type>
<position>208.5,-65.5</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>433 </input>
<output>
<ID>OUT</ID>425 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>502</ID>
<type>AI_XOR2</type>
<position>201.5,-65.5</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>434 </input>
<output>
<ID>OUT</ID>426 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>503</ID>
<type>DA_FROM</type>
<position>195.5,-60.5</position>
<input>
<ID>IN_0</ID>430 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>504</ID>
<type>DA_FROM</type>
<position>189,-60</position>
<input>
<ID>IN_0</ID>429 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>505</ID>
<type>DA_FROM</type>
<position>184,-60</position>
<input>
<ID>IN_0</ID>428 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>506</ID>
<type>DA_FROM</type>
<position>177.5,-59.5</position>
<input>
<ID>IN_0</ID>427 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>507</ID>
<type>AI_XOR2</type>
<position>196.5,-66.5</position>
<input>
<ID>IN_0</ID>444 </input>
<input>
<ID>IN_1</ID>430 </input>
<output>
<ID>OUT</ID>435 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>508</ID>
<type>AI_XOR2</type>
<position>190,-66.5</position>
<input>
<ID>IN_0</ID>444 </input>
<input>
<ID>IN_1</ID>429 </input>
<output>
<ID>OUT</ID>437 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>509</ID>
<type>AI_XOR2</type>
<position>185,-66.5</position>
<input>
<ID>IN_0</ID>444 </input>
<input>
<ID>IN_1</ID>428 </input>
<output>
<ID>OUT</ID>441 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>510</ID>
<type>AI_XOR2</type>
<position>178.5,-66.5</position>
<input>
<ID>IN_0</ID>444 </input>
<input>
<ID>IN_1</ID>427 </input>
<output>
<ID>OUT</ID>442 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>511</ID>
<type>AA_REGISTER4</type>
<position>194,-42.5</position>
<input>
<ID>IN_0</ID>458 </input>
<input>
<ID>IN_1</ID>457 </input>
<input>
<ID>IN_2</ID>456 </input>
<input>
<ID>IN_3</ID>455 </input>
<output>
<ID>OUT_0</ID>431 </output>
<output>
<ID>OUT_1</ID>432 </output>
<output>
<ID>OUT_2</ID>433 </output>
<output>
<ID>OUT_3</ID>434 </output>
<input>
<ID>clear</ID>468 </input>
<input>
<ID>clock</ID>467 </input>
<input>
<ID>count_enable</ID>469 </input>
<input>
<ID>count_up</ID>469 </input>
<input>
<ID>load</ID>470 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>512</ID>
<type>AA_AND2</type>
<position>197.5,-75</position>
<input>
<ID>IN_0</ID>443 </input>
<input>
<ID>IN_1</ID>435 </input>
<output>
<ID>OUT</ID>436 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>513</ID>
<type>AA_AND2</type>
<position>191,-75.5</position>
<input>
<ID>IN_0</ID>443 </input>
<input>
<ID>IN_1</ID>437 </input>
<output>
<ID>OUT</ID>438 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>514</ID>
<type>AA_AND2</type>
<position>186,-75.5</position>
<input>
<ID>IN_0</ID>443 </input>
<input>
<ID>IN_1</ID>441 </input>
<output>
<ID>OUT</ID>439 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>515</ID>
<type>AA_AND2</type>
<position>179.5,-75.5</position>
<input>
<ID>IN_0</ID>443 </input>
<input>
<ID>IN_1</ID>442 </input>
<output>
<ID>OUT</ID>440 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>516</ID>
<type>AE_SMALL_INVERTER</type>
<position>175,-71</position>
<input>
<ID>IN_0</ID>471 </input>
<output>
<ID>OUT_0</ID>443 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>519</ID>
<type>AA_AND4</type>
<position>-56.5,-26.5</position>
<input>
<ID>IN_0</ID>624 </input>
<input>
<ID>IN_1</ID>625 </input>
<input>
<ID>IN_2</ID>626 </input>
<input>
<ID>IN_3</ID>627 </input>
<output>
<ID>OUT</ID>630 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>521</ID>
<type>DA_FROM</type>
<position>201,-34.5</position>
<input>
<ID>IN_0</ID>470 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LD Acc</lparam></gate>
<gate>
<ID>522</ID>
<type>DA_FROM</type>
<position>166,-71</position>
<input>
<ID>IN_0</ID>471 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZero</lparam></gate>
<gate>
<ID>523</ID>
<type>DE_TO</type>
<position>148,-95.5</position>
<input>
<ID>IN_0</ID>446 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A4</lparam></gate>
<gate>
<ID>524</ID>
<type>DE_TO</type>
<position>142.5,-94</position>
<input>
<ID>IN_0</ID>447 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A5</lparam></gate>
<gate>
<ID>525</ID>
<type>DE_TO</type>
<position>149,-92.5</position>
<input>
<ID>IN_0</ID>448 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A6</lparam></gate>
<gate>
<ID>526</ID>
<type>DE_TO</type>
<position>143,-91</position>
<input>
<ID>IN_0</ID>449 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A7</lparam></gate>
<gate>
<ID>527</ID>
<type>BE_NOR4</type>
<position>155,-82</position>
<input>
<ID>IN_0</ID>449 </input>
<input>
<ID>IN_1</ID>448 </input>
<input>
<ID>IN_2</ID>447 </input>
<input>
<ID>IN_3</ID>446 </input>
<output>
<ID>OUT</ID>472 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>528</ID>
<type>DE_TO</type>
<position>155,-71</position>
<input>
<ID>IN_0</ID>472 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z7-4</lparam></gate>
<gate>
<ID>529</ID>
<type>AA_MUX_2x1</type>
<position>-56.5,-19.5</position>
<input>
<ID>IN_0</ID>315 </input>
<input>
<ID>IN_1</ID>630 </input>
<output>
<ID>OUT</ID>629 </output>
<input>
<ID>SEL_0</ID>631 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>531</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>271,-42</position>
<input>
<ID>ENABLE_0</ID>450 </input>
<input>
<ID>IN_0</ID>512 </input>
<input>
<ID>IN_1</ID>511 </input>
<input>
<ID>IN_2</ID>510 </input>
<input>
<ID>IN_3</ID>509 </input>
<output>
<ID>OUT_0</ID>508 </output>
<output>
<ID>OUT_1</ID>507 </output>
<output>
<ID>OUT_2</ID>506 </output>
<output>
<ID>OUT_3</ID>505 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>532</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>274.5,-32.5</position>
<input>
<ID>ENABLE_0</ID>395 </input>
<input>
<ID>IN_0</ID>516 </input>
<input>
<ID>IN_1</ID>515 </input>
<input>
<ID>IN_2</ID>514 </input>
<input>
<ID>IN_3</ID>513 </input>
<output>
<ID>OUT_0</ID>505 </output>
<output>
<ID>OUT_1</ID>506 </output>
<output>
<ID>OUT_2</ID>507 </output>
<output>
<ID>OUT_3</ID>508 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>533</ID>
<type>DA_FROM</type>
<position>264,-40.5</position>
<input>
<ID>IN_0</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>534</ID>
<type>DA_FROM</type>
<position>259.5,-41.5</position>
<input>
<ID>IN_0</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>535</ID>
<type>DA_FROM</type>
<position>254,-42.5</position>
<input>
<ID>IN_0</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>536</ID>
<type>DA_FROM</type>
<position>248,-43.5</position>
<input>
<ID>IN_0</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>537</ID>
<type>DA_FROM</type>
<position>323.5,-23.5</position>
<input>
<ID>IN_0</ID>513 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>538</ID>
<type>DA_FROM</type>
<position>319.5,-23</position>
<input>
<ID>IN_0</ID>514 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>539</ID>
<type>DA_FROM</type>
<position>316.5,-23</position>
<input>
<ID>IN_0</ID>515 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>540</ID>
<type>DA_FROM</type>
<position>313,-22.5</position>
<input>
<ID>IN_0</ID>516 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>541</ID>
<type>DA_FROM</type>
<position>275.5,-48</position>
<input>
<ID>IN_0</ID>517 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>542</ID>
<type>FF_GND</type>
<position>283,-47.5</position>
<output>
<ID>OUT_0</ID>518 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>543</ID>
<type>FF_GND</type>
<position>282,-35</position>
<output>
<ID>OUT_0</ID>519 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>544</ID>
<type>AE_FULLADDER_4BIT</type>
<position>287.5,-87</position>
<input>
<ID>IN_0</ID>486 </input>
<input>
<ID>IN_1</ID>488 </input>
<input>
<ID>IN_2</ID>489 </input>
<input>
<ID>IN_3</ID>490 </input>
<input>
<ID>IN_B_0</ID>473 </input>
<input>
<ID>IN_B_1</ID>474 </input>
<input>
<ID>IN_B_2</ID>475 </input>
<input>
<ID>IN_B_3</ID>476 </input>
<output>
<ID>OUT_0</ID>496 </output>
<output>
<ID>OUT_1</ID>497 </output>
<output>
<ID>OUT_2</ID>498 </output>
<output>
<ID>OUT_3</ID>499 </output>
<input>
<ID>carry_in</ID>500 </input>
<output>
<ID>carry_out</ID>524 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>545</ID>
<type>AI_XOR2</type>
<position>308.5,-65.5</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>481 </input>
<output>
<ID>OUT</ID>473 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>546</ID>
<type>AI_XOR2</type>
<position>302,-65.5</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>482 </input>
<output>
<ID>OUT</ID>474 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>547</ID>
<type>AI_XOR2</type>
<position>296.5,-65.5</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>483 </input>
<output>
<ID>OUT</ID>475 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>548</ID>
<type>AI_XOR2</type>
<position>289.5,-65.5</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>484 </input>
<output>
<ID>OUT</ID>476 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>549</ID>
<type>DA_FROM</type>
<position>283.5,-58.5</position>
<input>
<ID>IN_0</ID>480 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>550</ID>
<type>DA_FROM</type>
<position>277,-58</position>
<input>
<ID>IN_0</ID>479 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>551</ID>
<type>DA_FROM</type>
<position>272,-57.5</position>
<input>
<ID>IN_0</ID>478 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>552</ID>
<type>DA_FROM</type>
<position>265.5,-57.5</position>
<input>
<ID>IN_0</ID>477 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>553</ID>
<type>AI_XOR2</type>
<position>284.5,-66.5</position>
<input>
<ID>IN_0</ID>494 </input>
<input>
<ID>IN_1</ID>480 </input>
<output>
<ID>OUT</ID>485 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>554</ID>
<type>AI_XOR2</type>
<position>278,-66.5</position>
<input>
<ID>IN_0</ID>494 </input>
<input>
<ID>IN_1</ID>479 </input>
<output>
<ID>OUT</ID>487 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>555</ID>
<type>AI_XOR2</type>
<position>273,-66.5</position>
<input>
<ID>IN_0</ID>494 </input>
<input>
<ID>IN_1</ID>478 </input>
<output>
<ID>OUT</ID>491 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>556</ID>
<type>AI_XOR2</type>
<position>266.5,-66.5</position>
<input>
<ID>IN_0</ID>494 </input>
<input>
<ID>IN_1</ID>477 </input>
<output>
<ID>OUT</ID>492 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>557</ID>
<type>AA_REGISTER4</type>
<position>282,-42.5</position>
<input>
<ID>IN_0</ID>508 </input>
<input>
<ID>IN_1</ID>507 </input>
<input>
<ID>IN_2</ID>506 </input>
<input>
<ID>IN_3</ID>505 </input>
<output>
<ID>OUT_0</ID>481 </output>
<output>
<ID>OUT_1</ID>482 </output>
<output>
<ID>OUT_2</ID>483 </output>
<output>
<ID>OUT_3</ID>484 </output>
<input>
<ID>clear</ID>518 </input>
<input>
<ID>clock</ID>517 </input>
<input>
<ID>count_enable</ID>519 </input>
<input>
<ID>count_up</ID>519 </input>
<input>
<ID>load</ID>520 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>558</ID>
<type>AA_AND2</type>
<position>285.5,-75</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>485 </input>
<output>
<ID>OUT</ID>486 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>559</ID>
<type>AA_AND2</type>
<position>279,-75.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>487 </input>
<output>
<ID>OUT</ID>488 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>560</ID>
<type>AA_AND2</type>
<position>274,-75.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>491 </input>
<output>
<ID>OUT</ID>489 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>561</ID>
<type>AA_AND2</type>
<position>267.5,-75.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>490 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>562</ID>
<type>AE_SMALL_INVERTER</type>
<position>263,-71</position>
<input>
<ID>IN_0</ID>521 </input>
<output>
<ID>OUT_0</ID>493 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>563</ID>
<type>DA_FROM</type>
<position>-65,-19.5</position>
<input>
<ID>IN_0</ID>631 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID StatEn</lparam></gate>
<gate>
<ID>564</ID>
<type>AE_OR2</type>
<position>317.5,-65</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>494 </input>
<output>
<ID>OUT</ID>500 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>565</ID>
<type>AA_MUX_2x1</type>
<position>-58.5,-68.5</position>
<input>
<ID>IN_0</ID>303 </input>
<input>
<ID>IN_1</ID>336 </input>
<output>
<ID>OUT</ID>662 </output>
<input>
<ID>SEL_0</ID>632 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>566</ID>
<type>DA_FROM</type>
<position>-67,-68.5</position>
<input>
<ID>IN_0</ID>632 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID StatEn</lparam></gate>
<gate>
<ID>567</ID>
<type>DA_FROM</type>
<position>292,-33</position>
<input>
<ID>IN_0</ID>520 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LD Acc</lparam></gate>
<gate>
<ID>568</ID>
<type>DA_FROM</type>
<position>254,-71</position>
<input>
<ID>IN_0</ID>521 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZero</lparam></gate>
<gate>
<ID>569</ID>
<type>DE_TO</type>
<position>236,-95.5</position>
<input>
<ID>IN_0</ID>496 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>570</ID>
<type>DE_TO</type>
<position>230.5,-94</position>
<input>
<ID>IN_0</ID>497 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>571</ID>
<type>DE_TO</type>
<position>237,-92.5</position>
<input>
<ID>IN_0</ID>498 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>572</ID>
<type>DE_TO</type>
<position>231,-91</position>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>573</ID>
<type>BE_NOR4</type>
<position>243,-82</position>
<input>
<ID>IN_0</ID>499 </input>
<input>
<ID>IN_1</ID>498 </input>
<input>
<ID>IN_2</ID>497 </input>
<input>
<ID>IN_3</ID>496 </input>
<output>
<ID>OUT</ID>522 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>574</ID>
<type>DE_TO</type>
<position>243,-71</position>
<input>
<ID>IN_0</ID>522 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z3-0</lparam></gate>
<gate>
<ID>575</ID>
<type>AA_MUX_2x1</type>
<position>-44,-83.5</position>
<input>
<ID>IN_0</ID>294 </input>
<input>
<ID>IN_1</ID>692 </input>
<output>
<ID>OUT</ID>669 </output>
<input>
<ID>SEL_0</ID>668 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>576</ID>
<type>DA_FROM</type>
<position>-56,-83.5</position>
<input>
<ID>IN_0</ID>668 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID StatEn</lparam></gate>
<gate>
<ID>577</ID>
<type>AA_MUX_2x1</type>
<position>-22.5,-82.5</position>
<input>
<ID>IN_0</ID>298 </input>
<input>
<ID>IN_1</ID>704 </input>
<output>
<ID>OUT</ID>703 </output>
<input>
<ID>SEL_0</ID>702 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>578</ID>
<type>DA_FROM</type>
<position>-32.5,-68.5</position>
<input>
<ID>IN_0</ID>702 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID StatEn</lparam></gate>
<gate>
<ID>586</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>311,-42</position>
<input>
<ID>ENABLE_0</ID>531 </input>
<input>
<ID>IN_0</ID>481 </input>
<input>
<ID>IN_1</ID>482 </input>
<input>
<ID>IN_2</ID>483 </input>
<input>
<ID>IN_3</ID>484 </input>
<output>
<ID>OUT_0</ID>513 </output>
<output>
<ID>OUT_1</ID>514 </output>
<output>
<ID>OUT_2</ID>515 </output>
<output>
<ID>OUT_3</ID>516 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>588</ID>
<type>DA_FROM</type>
<position>307,-38</position>
<input>
<ID>IN_0</ID>531 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Acc-Bus</lparam></gate>
<gate>
<ID>589</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>222.5,-42</position>
<input>
<ID>ENABLE_0</ID>532 </input>
<input>
<ID>IN_0</ID>431 </input>
<input>
<ID>IN_1</ID>432 </input>
<input>
<ID>IN_2</ID>433 </input>
<input>
<ID>IN_3</ID>434 </input>
<output>
<ID>OUT_0</ID>463 </output>
<output>
<ID>OUT_1</ID>464 </output>
<output>
<ID>OUT_2</ID>465 </output>
<output>
<ID>OUT_3</ID>466 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>590</ID>
<type>DA_FROM</type>
<position>218.5,-37.5</position>
<input>
<ID>IN_0</ID>532 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Acc-Bus</lparam></gate>
<gate>
<ID>591</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>133.5,-42</position>
<input>
<ID>ENABLE_0</ID>533 </input>
<input>
<ID>IN_0</ID>375 </input>
<input>
<ID>IN_1</ID>376 </input>
<input>
<ID>IN_2</ID>377 </input>
<input>
<ID>IN_3</ID>378 </input>
<output>
<ID>OUT_0</ID>407 </output>
<output>
<ID>OUT_1</ID>408 </output>
<output>
<ID>OUT_2</ID>409 </output>
<output>
<ID>OUT_3</ID>410 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>592</ID>
<type>DA_FROM</type>
<position>131,-37.5</position>
<input>
<ID>IN_0</ID>533 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Acc-Bus</lparam></gate>
<gate>
<ID>593</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>42,-43</position>
<input>
<ID>ENABLE_0</ID>534 </input>
<input>
<ID>IN_0</ID>317 </input>
<input>
<ID>IN_1</ID>318 </input>
<input>
<ID>IN_2</ID>319 </input>
<input>
<ID>IN_3</ID>320 </input>
<output>
<ID>OUT_0</ID>351 </output>
<output>
<ID>OUT_1</ID>352 </output>
<output>
<ID>OUT_2</ID>353 </output>
<output>
<ID>OUT_3</ID>354 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>594</ID>
<type>DA_FROM</type>
<position>39.5,-38.5</position>
<input>
<ID>IN_0</ID>534 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Acc-Bus</lparam></gate>
<gate>
<ID>596</ID>
<type>DA_FROM</type>
<position>326,-59</position>
<input>
<ID>IN_0</ID>495 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBA</lparam></gate>
<gate>
<ID>597</ID>
<type>DA_FROM</type>
<position>324.5,-54.5</position>
<input>
<ID>IN_0</ID>494 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBB</lparam></gate>
<gate>
<ID>599</ID>
<type>DA_FROM</type>
<position>236.5,-58</position>
<input>
<ID>IN_0</ID>445 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBA</lparam></gate>
<gate>
<ID>600</ID>
<type>DA_FROM</type>
<position>235,-53.5</position>
<input>
<ID>IN_0</ID>444 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBB</lparam></gate>
<gate>
<ID>601</ID>
<type>DA_FROM</type>
<position>139.5,-58</position>
<input>
<ID>IN_0</ID>389 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBA</lparam></gate>
<gate>
<ID>602</ID>
<type>DA_FROM</type>
<position>138,-53.5</position>
<input>
<ID>IN_0</ID>388 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBB</lparam></gate>
<gate>
<ID>603</ID>
<type>DA_FROM</type>
<position>-52,-36.5</position>
<input>
<ID>IN_0</ID>626 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z7-4</lparam></gate>
<gate>
<ID>604</ID>
<type>DA_FROM</type>
<position>-49,-36.5</position>
<input>
<ID>IN_0</ID>627 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z3-0</lparam></gate>
<gate>
<ID>605</ID>
<type>DA_FROM</type>
<position>51,-55.5</position>
<input>
<ID>IN_0</ID>332 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBA</lparam></gate>
<gate>
<ID>606</ID>
<type>DA_FROM</type>
<position>49,-51.5</position>
<input>
<ID>IN_0</ID>331 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBB</lparam></gate>
<gate>
<ID>608</ID>
<type>DA_FROM</type>
<position>0,-37</position>
<input>
<ID>IN_0</ID>537 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD Acc</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_LABEL</type>
<position>61,-9</position>
<gparam>LABEL_TEXT Accumulator</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>660</ID>
<type>AA_TOGGLE</type>
<position>287,-6</position>
<output>
<ID>OUT_0</ID>719 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>335</ID>
<type>AE_FULLADDER_4BIT</type>
<position>19.5,-88</position>
<input>
<ID>IN_0</ID>322 </input>
<input>
<ID>IN_1</ID>324 </input>
<input>
<ID>IN_2</ID>325 </input>
<input>
<ID>IN_3</ID>326 </input>
<input>
<ID>IN_B_0</ID>287 </input>
<input>
<ID>IN_B_1</ID>288 </input>
<input>
<ID>IN_B_2</ID>289 </input>
<input>
<ID>IN_B_3</ID>290 </input>
<output>
<ID>OUT_0</ID>661 </output>
<output>
<ID>OUT_1</ID>334 </output>
<output>
<ID>OUT_2</ID>335 </output>
<output>
<ID>OUT_3</ID>336 </output>
<input>
<ID>carry_in</ID>414 </input>
<output>
<ID>carry_out</ID>692 </output>
<output>
<ID>overflow</ID>704 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>336</ID>
<type>AE_DFF_LOW</type>
<position>-41,-78</position>
<input>
<ID>IN_0</ID>669 </input>
<output>
<ID>OUT_0</ID>294 </output>
<input>
<ID>clear</ID>292 </input>
<input>
<ID>clock</ID>293 </input>
<input>
<ID>set</ID>291 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>337</ID>
<type>EE_VDD</type>
<position>-47,-78</position>
<output>
<ID>OUT_0</ID>291 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>338</ID>
<type>AI_XOR2</type>
<position>40.5,-66.5</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>317 </input>
<output>
<ID>OUT</ID>287 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>339</ID>
<type>AI_XOR2</type>
<position>34,-66.5</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>318 </input>
<output>
<ID>OUT</ID>288 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>340</ID>
<type>AI_XOR2</type>
<position>28.5,-66.5</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>319 </input>
<output>
<ID>OUT</ID>289 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>AI_XOR2</type>
<position>21.5,-66.5</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>320 </input>
<output>
<ID>OUT</ID>290 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>342</ID>
<type>EE_VDD</type>
<position>-31,-78</position>
<output>
<ID>OUT_0</ID>292 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>343</ID>
<type>DA_FROM</type>
<position>15.5,-61</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>344</ID>
<type>DA_FROM</type>
<position>9,-60</position>
<input>
<ID>IN_0</ID>309 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>345</ID>
<type>DA_FROM</type>
<position>4,-60.5</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>346</ID>
<type>DA_FROM</type>
<position>-2.5,-58.5</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>347</ID>
<type>GA_LED</type>
<position>-46.5,-89</position>
<input>
<ID>N_in1</ID>704 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>348</ID>
<type>DA_FROM</type>
<position>-40,-83.5</position>
<input>
<ID>IN_0</ID>293 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>349</ID>
<type>GA_LED</type>
<position>-43,-70.5</position>
<input>
<ID>N_in2</ID>294 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>350</ID>
<type>GA_LED</type>
<position>-50,-87</position>
<input>
<ID>N_in1</ID>692 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>351</ID>
<type>AI_XOR2</type>
<position>16.5,-67.5</position>
<input>
<ID>IN_0</ID>331 </input>
<input>
<ID>IN_1</ID>310 </input>
<output>
<ID>OUT</ID>321 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>352</ID>
<type>AI_XOR2</type>
<position>10,-67.5</position>
<input>
<ID>IN_0</ID>331 </input>
<input>
<ID>IN_1</ID>309 </input>
<output>
<ID>OUT</ID>323 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>353</ID>
<type>AI_XOR2</type>
<position>5,-67.5</position>
<input>
<ID>IN_0</ID>331 </input>
<input>
<ID>IN_1</ID>308 </input>
<output>
<ID>OUT</ID>327 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>354</ID>
<type>AI_XOR2</type>
<position>-1.5,-67.5</position>
<input>
<ID>IN_0</ID>331 </input>
<input>
<ID>IN_1</ID>307 </input>
<output>
<ID>OUT</ID>328 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>355</ID>
<type>DE_TO</type>
<position>-46,-73.5</position>
<input>
<ID>IN_0</ID>294 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Carry</lparam></gate>
<gate>
<ID>356</ID>
<type>AE_DFF_LOW</type>
<position>-20.5,-77.5</position>
<input>
<ID>IN_0</ID>703 </input>
<output>
<ID>OUT_0</ID>298 </output>
<input>
<ID>clear</ID>296 </input>
<input>
<ID>clock</ID>297 </input>
<input>
<ID>set</ID>295 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>357</ID>
<type>EE_VDD</type>
<position>-26.5,-77.5</position>
<output>
<ID>OUT_0</ID>295 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>358</ID>
<type>EE_VDD</type>
<position>-13,-77.5</position>
<output>
<ID>OUT_0</ID>296 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>359</ID>
<type>DA_FROM</type>
<position>-19.5,-83</position>
<input>
<ID>IN_0</ID>297 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>360</ID>
<type>GA_LED</type>
<position>-22.5,-70</position>
<input>
<ID>N_in2</ID>298 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>362</ID>
<type>DE_TO</type>
<position>-24.5,-72.5</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID oVerflow</lparam></gate>
<gate>
<ID>364</ID>
<type>AE_DFF_LOW</type>
<position>-52,-59</position>
<input>
<ID>IN_0</ID>662 </input>
<output>
<ID>OUT_0</ID>303 </output>
<input>
<ID>clear</ID>301 </input>
<input>
<ID>clock</ID>302 </input>
<input>
<ID>set</ID>299 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>366</ID>
<type>EE_VDD</type>
<position>-58,-59</position>
<output>
<ID>OUT_0</ID>299 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>368</ID>
<type>EE_VDD</type>
<position>-46,-59</position>
<output>
<ID>OUT_0</ID>301 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_REGISTER4</type>
<position>14,-43.5</position>
<input>
<ID>IN_0</ID>346 </input>
<input>
<ID>IN_1</ID>345 </input>
<input>
<ID>IN_2</ID>344 </input>
<input>
<ID>IN_3</ID>343 </input>
<output>
<ID>OUT_0</ID>317 </output>
<output>
<ID>OUT_1</ID>318 </output>
<output>
<ID>OUT_2</ID>319 </output>
<output>
<ID>OUT_3</ID>320 </output>
<input>
<ID>clear</ID>356 </input>
<input>
<ID>clock</ID>355 </input>
<input>
<ID>count_enable</ID>357 </input>
<input>
<ID>count_up</ID>357 </input>
<input>
<ID>load</ID>537 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>370</ID>
<type>DA_FROM</type>
<position>-51,-64.5</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>371</ID>
<type>AA_AND2</type>
<position>17.5,-76</position>
<input>
<ID>IN_0</ID>329 </input>
<input>
<ID>IN_1</ID>321 </input>
<output>
<ID>OUT</ID>322 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>372</ID>
<type>AA_AND2</type>
<position>11,-76.5</position>
<input>
<ID>IN_0</ID>329 </input>
<input>
<ID>IN_1</ID>323 </input>
<output>
<ID>OUT</ID>324 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>373</ID>
<type>AA_AND2</type>
<position>6,-76.5</position>
<input>
<ID>IN_0</ID>329 </input>
<input>
<ID>IN_1</ID>327 </input>
<output>
<ID>OUT</ID>325 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>374</ID>
<type>AA_AND2</type>
<position>-0.5,-76.5</position>
<input>
<ID>IN_0</ID>329 </input>
<input>
<ID>IN_1</ID>328 </input>
<output>
<ID>OUT</ID>326 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>375</ID>
<type>GA_LED</type>
<position>-54,-51.5</position>
<input>
<ID>N_in2</ID>303 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>376</ID>
<type>AE_SMALL_INVERTER</type>
<position>-5,-72</position>
<input>
<ID>IN_0</ID>417 </input>
<output>
<ID>OUT_0</ID>329 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>377</ID>
<type>DE_TO</type>
<position>-57,-54.5</position>
<input>
<ID>IN_0</ID>303 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID sigN</lparam></gate>
<gate>
<ID>379</ID>
<type>AE_DFF_LOW</type>
<position>-54.5,-13</position>
<input>
<ID>IN_0</ID>629 </input>
<output>
<ID>OUT_0</ID>315 </output>
<input>
<ID>clear</ID>306 </input>
<input>
<ID>clock</ID>311 </input>
<input>
<ID>set</ID>304 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>381</ID>
<type>EE_VDD</type>
<position>-58.5,-12</position>
<output>
<ID>OUT_0</ID>304 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>382</ID>
<type>DA_FROM</type>
<position>18,-33.5</position>
<input>
<ID>IN_0</ID>369 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus-Acc</lparam></gate>
<gate>
<ID>383</ID>
<type>EE_VDD</type>
<position>-46.5,-12</position>
<output>
<ID>OUT_0</ID>306 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>384</ID>
<type>DA_FROM</type>
<position>102,-32.5</position>
<input>
<ID>IN_0</ID>370 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus-Acc</lparam></gate>
<gate>
<ID>385</ID>
<type>DA_FROM</type>
<position>191.5,-32.5</position>
<input>
<ID>IN_0</ID>394 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus-Acc</lparam></gate>
<gate>
<ID>386</ID>
<type>DA_FROM</type>
<position>281,-31.5</position>
<input>
<ID>IN_0</ID>395 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus-Acc</lparam></gate>
<gate>
<ID>387</ID>
<type>DA_FROM</type>
<position>3,-29.5</position>
<input>
<ID>IN_0</ID>396 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Res-Acc</lparam></gate>
<gate>
<ID>388</ID>
<type>DA_FROM</type>
<position>-52,-19.5</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-62.5,113,-51.5</points>
<connection>
<GID>435</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113,-51.5,132,-51.5</points>
<intersection>113 0</intersection>
<intersection>120 3</intersection>
<intersection>125.5 7</intersection>
<intersection>132 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>120,-62.5,120,-51.5</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>132,-62.5,132,-51.5</points>
<connection>
<GID>432</GID>
<name>IN_0</name></connection>
<intersection>-58 10</intersection>
<intersection>-51.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>125.5,-62.5,125.5,-51.5</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>132,-58,137.5,-58</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<intersection>132 6</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-95.5,111.5,-91</points>
<connection>
<GID>431</GID>
<name>OUT_0</name></connection>
<intersection>-95.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>60.5,-95.5,111.5,-95.5</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>68.5 8</intersection>
<intersection>111.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>68.5,-95.5,68.5,-85</points>
<connection>
<GID>480</GID>
<name>IN_3</name></connection>
<intersection>-95.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-94,110.5,-91</points>
<connection>
<GID>431</GID>
<name>OUT_1</name></connection>
<intersection>-94 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>55,-94,110.5,-94</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<intersection>66.5 8</intersection>
<intersection>110.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>66.5,-94,66.5,-85</points>
<connection>
<GID>480</GID>
<name>IN_2</name></connection>
<intersection>-94 7</intersection></vsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-92.5,109.5,-91</points>
<connection>
<GID>431</GID>
<name>OUT_2</name></connection>
<intersection>-92.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>61.5,-92.5,109.5,-92.5</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<intersection>64.5 8</intersection>
<intersection>109.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>64.5,-92.5,64.5,-85</points>
<connection>
<GID>480</GID>
<name>IN_1</name></connection>
<intersection>-92.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>55.5,-91,108.5,-91</points>
<connection>
<GID>431</GID>
<name>OUT_3</name></connection>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>62.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>62.5,-91,62.5,-85</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>-91 7</intersection></vsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,-32.5,189.5,-32.5</points>
<connection>
<GID>486</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>385</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-32.5,278,-31.5</points>
<intersection>-32.5 1</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277.5,-32.5,278,-32.5</points>
<connection>
<GID>532</GID>
<name>ENABLE_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>278,-31.5,279,-31.5</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-40,3,-31.5</points>
<connection>
<GID>395</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>387</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-39,93.5,-24.5</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<connection>
<GID>418</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-39,183,-31</points>
<connection>
<GID>485</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>410</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95.5,-40.5,100.5,-40.5</points>
<connection>
<GID>418</GID>
<name>OUT_3</name></connection>
<connection>
<GID>450</GID>
<name>IN_3</name></connection>
<intersection>95.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>95.5,-40.5,95.5,-34.5</points>
<connection>
<GID>419</GID>
<name>OUT_0</name></connection>
<intersection>-40.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95.5,-41.5,100.5,-41.5</points>
<connection>
<GID>418</GID>
<name>OUT_2</name></connection>
<connection>
<GID>450</GID>
<name>IN_2</name></connection>
<intersection>96.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>96.5,-41.5,96.5,-34.5</points>
<connection>
<GID>419</GID>
<name>OUT_1</name></connection>
<intersection>-41.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95.5,-42.5,100.5,-42.5</points>
<connection>
<GID>418</GID>
<name>OUT_1</name></connection>
<connection>
<GID>450</GID>
<name>IN_1</name></connection>
<intersection>97.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>97.5,-42.5,97.5,-34.5</points>
<connection>
<GID>419</GID>
<name>OUT_2</name></connection>
<intersection>-42.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95.5,-43.5,100.5,-43.5</points>
<connection>
<GID>418</GID>
<name>OUT_0</name></connection>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>98.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>98.5,-43.5,98.5,-34.5</points>
<connection>
<GID>419</GID>
<name>OUT_3</name></connection>
<intersection>-43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88.5,-40.5,91.5,-40.5</points>
<connection>
<GID>418</GID>
<name>IN_3</name></connection>
<connection>
<GID>420</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>84,-41.5,91.5,-41.5</points>
<connection>
<GID>418</GID>
<name>IN_2</name></connection>
<connection>
<GID>421</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78.5,-42.5,91.5,-42.5</points>
<connection>
<GID>418</GID>
<name>IN_1</name></connection>
<connection>
<GID>422</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72.5,-43.5,91.5,-43.5</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<connection>
<GID>423</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-30.5,98.5,-30</points>
<connection>
<GID>419</GID>
<name>IN_3</name></connection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>98.5,-30,148,-30</points>
<intersection>98.5 0</intersection>
<intersection>148 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>148,-43.5,148,-24.5</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>-43.5 5</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>135.5,-43.5,148,-43.5</points>
<connection>
<GID>591</GID>
<name>OUT_0</name></connection>
<intersection>148 3</intersection></hsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-42.5,144,-24</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<intersection>-42.5 10</intersection>
<intersection>-29 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>97.5,-29,144,-29</points>
<intersection>97.5 8</intersection>
<intersection>144 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>97.5,-30.5,97.5,-29</points>
<connection>
<GID>419</GID>
<name>IN_2</name></connection>
<intersection>-29 7</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>135.5,-42.5,144,-42.5</points>
<connection>
<GID>591</GID>
<name>OUT_1</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-30.5,96.5,-27.5</points>
<connection>
<GID>419</GID>
<name>IN_1</name></connection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>96.5,-27.5,140,-27.5</points>
<intersection>96.5 0</intersection>
<intersection>140 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>140,-41.5,140,-23.5</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<intersection>-41.5 9</intersection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>135.5,-41.5,140,-41.5</points>
<connection>
<GID>591</GID>
<name>OUT_2</name></connection>
<intersection>140 7</intersection></hsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-30.5,95.5,-26</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>-26 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>137,-40.5,137,-23.5</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>-40.5 4</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-26,137,-26</points>
<intersection>95.5 0</intersection>
<intersection>137 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>135.5,-40.5,137,-40.5</points>
<connection>
<GID>591</GID>
<name>OUT_3</name></connection>
<intersection>137 1</intersection></hsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-48,103.5,-46.5</points>
<connection>
<GID>450</GID>
<name>clock</name></connection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-48,103.5,-48</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-46.5,105.5,-46.5</points>
<connection>
<GID>429</GID>
<name>OUT_0</name></connection>
<connection>
<GID>450</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-37.5,104.5,-36</points>
<connection>
<GID>430</GID>
<name>OUT_0</name></connection>
<connection>
<GID>450</GID>
<name>count_enable</name></connection>
<intersection>-37.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-37.5,105.5,-37.5</points>
<connection>
<GID>450</GID>
<name>count_up</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-86,102,-86</points>
<connection>
<GID>431</GID>
<name>carry_out</name></connection>
<intersection>27.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>27.5,-87,27.5,-86</points>
<connection>
<GID>335</GID>
<name>carry_in</name></connection>
<intersection>-86 1</intersection></vsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-37.5,103.5,-33.5</points>
<connection>
<GID>450</GID>
<name>load</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-33.5,112.5,-33.5</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<intersection>103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78.5,-71,83.5,-71</points>
<connection>
<GID>455</GID>
<name>IN_0</name></connection>
<connection>
<GID>464</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-68.5,-7,-68.5</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>-7 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-7,-72,-7,-68.5</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>-68.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31.5,-79.5,-31.5,-63</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<connection>
<GID>397</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-78,65.5,-73</points>
<connection>
<GID>480</GID>
<name>OUT</name></connection>
<connection>
<GID>482</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220.5,-83,220.5,-68.5</points>
<connection>
<GID>499</GID>
<name>OUT</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>204.5,-83,220.5,-83</points>
<connection>
<GID>498</GID>
<name>IN_B_0</name></connection>
<intersection>220.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214,-82,214,-68.5</points>
<connection>
<GID>500</GID>
<name>OUT</name></connection>
<intersection>-82 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>203.5,-82,214,-82</points>
<intersection>203.5 4</intersection>
<intersection>214 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>203.5,-83,203.5,-82</points>
<connection>
<GID>498</GID>
<name>IN_B_1</name></connection>
<intersection>-82 3</intersection></vsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202.5,-83,202.5,-81</points>
<connection>
<GID>498</GID>
<name>IN_B_2</name></connection>
<intersection>-81 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>208.5,-81,208.5,-68.5</points>
<connection>
<GID>501</GID>
<name>OUT</name></connection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>202.5,-81,208.5,-81</points>
<intersection>202.5 0</intersection>
<intersection>208.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,-83,201.5,-68.5</points>
<connection>
<GID>502</GID>
<name>OUT</name></connection>
<connection>
<GID>498</GID>
<name>IN_B_3</name></connection></vsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177.5,-63.5,177.5,-61.5</points>
<connection>
<GID>510</GID>
<name>IN_1</name></connection>
<connection>
<GID>506</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-63.5,184,-62</points>
<connection>
<GID>509</GID>
<name>IN_1</name></connection>
<connection>
<GID>505</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-63.5,189,-62</points>
<connection>
<GID>508</GID>
<name>IN_1</name></connection>
<connection>
<GID>504</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>195.5,-63.5,195.5,-62.5</points>
<connection>
<GID>507</GID>
<name>IN_1</name></connection>
<connection>
<GID>503</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-62.5,219.5,-43.5</points>
<connection>
<GID>499</GID>
<name>IN_1</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198,-43.5,220.5,-43.5</points>
<connection>
<GID>511</GID>
<name>OUT_0</name></connection>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<intersection>219.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-62.5,213,-42.5</points>
<connection>
<GID>500</GID>
<name>IN_1</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198,-42.5,220.5,-42.5</points>
<connection>
<GID>511</GID>
<name>OUT_1</name></connection>
<connection>
<GID>589</GID>
<name>IN_1</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-62.5,207.5,-41.5</points>
<connection>
<GID>501</GID>
<name>IN_1</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198,-41.5,220.5,-41.5</points>
<connection>
<GID>511</GID>
<name>OUT_2</name></connection>
<connection>
<GID>589</GID>
<name>IN_2</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200.5,-62.5,200.5,-40.5</points>
<connection>
<GID>502</GID>
<name>IN_1</name></connection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198,-40.5,220.5,-40.5</points>
<connection>
<GID>511</GID>
<name>OUT_3</name></connection>
<connection>
<GID>589</GID>
<name>IN_3</name></connection>
<intersection>200.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,-72,196.5,-69.5</points>
<connection>
<GID>512</GID>
<name>IN_1</name></connection>
<connection>
<GID>507</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-83,197.5,-78</points>
<connection>
<GID>512</GID>
<name>OUT</name></connection>
<connection>
<GID>498</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-72.5,190,-69.5</points>
<connection>
<GID>513</GID>
<name>IN_1</name></connection>
<connection>
<GID>508</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,-83,196.5,-79.5</points>
<connection>
<GID>498</GID>
<name>IN_1</name></connection>
<intersection>-79.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>191,-79.5,196.5,-79.5</points>
<intersection>191 3</intersection>
<intersection>196.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>191,-79.5,191,-78.5</points>
<connection>
<GID>513</GID>
<name>OUT</name></connection>
<intersection>-79.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,-83,195.5,-80.5</points>
<connection>
<GID>498</GID>
<name>IN_2</name></connection>
<intersection>-80.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>186,-80.5,186,-78.5</points>
<connection>
<GID>514</GID>
<name>OUT</name></connection>
<intersection>-80.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>186,-80.5,195.5,-80.5</points>
<intersection>186 1</intersection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-83,194.5,-81.5</points>
<connection>
<GID>498</GID>
<name>IN_3</name></connection>
<intersection>-81.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>179.5,-81.5,179.5,-78.5</points>
<connection>
<GID>515</GID>
<name>OUT</name></connection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>179.5,-81.5,194.5,-81.5</points>
<intersection>179.5 1</intersection>
<intersection>194.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-72.5,185,-69.5</points>
<connection>
<GID>514</GID>
<name>IN_1</name></connection>
<connection>
<GID>509</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-72.5,178.5,-69.5</points>
<connection>
<GID>515</GID>
<name>IN_1</name></connection>
<connection>
<GID>510</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180.5,-72.5,180.5,-71</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177,-71,198.5,-71</points>
<connection>
<GID>516</GID>
<name>OUT_0</name></connection>
<intersection>180.5 0</intersection>
<intersection>187 3</intersection>
<intersection>192 5</intersection>
<intersection>198.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>187,-72.5,187,-71</points>
<connection>
<GID>514</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>192,-72.5,192,-71</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>198.5,-72,198.5,-71</points>
<connection>
<GID>512</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-63.5,179.5,-52.5</points>
<connection>
<GID>510</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>179.5,-52.5,197.5,-52.5</points>
<intersection>179.5 0</intersection>
<intersection>186 7</intersection>
<intersection>191 6</intersection>
<intersection>197.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>197.5,-63.5,197.5,-52.5</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>-53.5 10</intersection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>191,-63.5,191,-52.5</points>
<connection>
<GID>508</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>186,-63.5,186,-52.5</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>197.5,-53.5,233,-53.5</points>
<connection>
<GID>600</GID>
<name>IN_0</name></connection>
<intersection>197.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202.5,-62.5,202.5,-51.5</points>
<connection>
<GID>502</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,-51.5,221.5,-51.5</points>
<intersection>202.5 0</intersection>
<intersection>209.5 3</intersection>
<intersection>215 7</intersection>
<intersection>221.5 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>209.5,-62.5,209.5,-51.5</points>
<connection>
<GID>501</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>221.5,-62.5,221.5,-51.5</points>
<connection>
<GID>499</GID>
<name>IN_0</name></connection>
<intersection>-58 10</intersection>
<intersection>-51.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>215,-62.5,215,-51.5</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>221.5,-58,234.5,-58</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<intersection>221.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-95.5,201,-91</points>
<connection>
<GID>498</GID>
<name>OUT_0</name></connection>
<intersection>-95.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>150,-95.5,201,-95.5</points>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<intersection>158 8</intersection>
<intersection>201 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>158,-95.5,158,-85</points>
<connection>
<GID>527</GID>
<name>IN_3</name></connection>
<intersection>-95.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200,-94,200,-91</points>
<connection>
<GID>498</GID>
<name>OUT_1</name></connection>
<intersection>-94 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>144.5,-94,200,-94</points>
<connection>
<GID>524</GID>
<name>IN_0</name></connection>
<intersection>156 8</intersection>
<intersection>200 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>156,-94,156,-85</points>
<connection>
<GID>527</GID>
<name>IN_2</name></connection>
<intersection>-94 7</intersection></vsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-92.5,199,-91</points>
<connection>
<GID>498</GID>
<name>OUT_2</name></connection>
<intersection>-92.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>151,-92.5,199,-92.5</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<intersection>154 8</intersection>
<intersection>199 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>154,-92.5,154,-85</points>
<connection>
<GID>527</GID>
<name>IN_1</name></connection>
<intersection>-92.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>145,-91,198,-91</points>
<connection>
<GID>498</GID>
<name>OUT_3</name></connection>
<connection>
<GID>526</GID>
<name>IN_0</name></connection>
<intersection>152 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>152,-91,152,-85</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<intersection>-91 7</intersection></vsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-39,271,-29</points>
<connection>
<GID>531</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>411</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>185,-40.5,190,-40.5</points>
<connection>
<GID>485</GID>
<name>OUT_3</name></connection>
<connection>
<GID>511</GID>
<name>IN_3</name></connection>
<intersection>185 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>185,-40.5,185,-34.5</points>
<connection>
<GID>486</GID>
<name>OUT_0</name></connection>
<intersection>-40.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>185,-41.5,190,-41.5</points>
<connection>
<GID>485</GID>
<name>OUT_2</name></connection>
<connection>
<GID>511</GID>
<name>IN_2</name></connection>
<intersection>186 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>186,-41.5,186,-34.5</points>
<connection>
<GID>486</GID>
<name>OUT_1</name></connection>
<intersection>-41.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>185,-42.5,190,-42.5</points>
<connection>
<GID>485</GID>
<name>OUT_1</name></connection>
<connection>
<GID>511</GID>
<name>IN_1</name></connection>
<intersection>187 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>187,-42.5,187,-34.5</points>
<connection>
<GID>486</GID>
<name>OUT_2</name></connection>
<intersection>-42.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>185,-43.5,190,-43.5</points>
<connection>
<GID>485</GID>
<name>OUT_0</name></connection>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>188 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>188,-43.5,188,-34.5</points>
<connection>
<GID>486</GID>
<name>OUT_3</name></connection>
<intersection>-43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>178,-40.5,181,-40.5</points>
<connection>
<GID>485</GID>
<name>IN_3</name></connection>
<connection>
<GID>487</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>173.5,-41.5,181,-41.5</points>
<connection>
<GID>485</GID>
<name>IN_2</name></connection>
<connection>
<GID>488</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>168,-42.5,181,-42.5</points>
<connection>
<GID>485</GID>
<name>IN_1</name></connection>
<connection>
<GID>489</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-43.5,181,-43.5</points>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,-30.5,188,-29.5</points>
<connection>
<GID>486</GID>
<name>IN_3</name></connection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>188,-29.5,235.5,-29.5</points>
<intersection>188 0</intersection>
<intersection>235.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>235.5,-43.5,235.5,-26.5</points>
<connection>
<GID>491</GID>
<name>IN_0</name></connection>
<intersection>-43.5 5</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>224.5,-43.5,235.5,-43.5</points>
<connection>
<GID>589</GID>
<name>OUT_0</name></connection>
<intersection>235.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-42.5,231.5,-26</points>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<intersection>-42.5 10</intersection>
<intersection>-28.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>187,-28.5,231.5,-28.5</points>
<intersection>187 8</intersection>
<intersection>231.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>187,-30.5,187,-28.5</points>
<connection>
<GID>486</GID>
<name>IN_2</name></connection>
<intersection>-28.5 7</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>224.5,-42.5,231.5,-42.5</points>
<connection>
<GID>589</GID>
<name>OUT_1</name></connection>
<intersection>231.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-30.5,186,-27.5</points>
<connection>
<GID>486</GID>
<name>IN_1</name></connection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>186,-27.5,227.5,-27.5</points>
<intersection>186 0</intersection>
<intersection>227.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>227.5,-41.5,227.5,-25.5</points>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<intersection>-41.5 9</intersection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>224.5,-41.5,227.5,-41.5</points>
<connection>
<GID>589</GID>
<name>OUT_2</name></connection>
<intersection>227.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-30.5,185,-26.5</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>-26.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>224.5,-40.5,224.5,-25.5</points>
<connection>
<GID>589</GID>
<name>OUT_3</name></connection>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>185,-26.5,224.5,-26.5</points>
<intersection>185 0</intersection>
<intersection>224.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193,-48,193,-46.5</points>
<connection>
<GID>511</GID>
<name>clock</name></connection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,-48,193,-48</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-46.5,195,-46.5</points>
<connection>
<GID>496</GID>
<name>OUT_0</name></connection>
<connection>
<GID>511</GID>
<name>clear</name></connection></hsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>194,-37.5,195,-37.5</points>
<connection>
<GID>511</GID>
<name>count_up</name></connection>
<connection>
<GID>511</GID>
<name>count_enable</name></connection>
<intersection>194 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>194,-37.5,194,-37</points>
<connection>
<GID>497</GID>
<name>OUT_0</name></connection>
<intersection>-37.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193,-37.5,193,-34.5</points>
<connection>
<GID>511</GID>
<name>load</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193,-34.5,199,-34.5</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>193 0</intersection></hsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>168,-71,173,-71</points>
<connection>
<GID>516</GID>
<name>IN_0</name></connection>
<connection>
<GID>522</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-78,155,-73</points>
<connection>
<GID>528</GID>
<name>IN_0</name></connection>
<connection>
<GID>527</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308.5,-83,308.5,-68.5</points>
<connection>
<GID>545</GID>
<name>OUT</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292.5,-83,308.5,-83</points>
<connection>
<GID>544</GID>
<name>IN_B_0</name></connection>
<intersection>308.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-82,302,-68.5</points>
<connection>
<GID>546</GID>
<name>OUT</name></connection>
<intersection>-82 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>291.5,-82,302,-82</points>
<intersection>291.5 4</intersection>
<intersection>302 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>291.5,-83,291.5,-82</points>
<connection>
<GID>544</GID>
<name>IN_B_1</name></connection>
<intersection>-82 3</intersection></vsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-83,290.5,-81</points>
<connection>
<GID>544</GID>
<name>IN_B_2</name></connection>
<intersection>-81 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>296.5,-81,296.5,-68.5</points>
<connection>
<GID>547</GID>
<name>OUT</name></connection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>290.5,-81,296.5,-81</points>
<intersection>290.5 0</intersection>
<intersection>296.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289.5,-83,289.5,-68.5</points>
<connection>
<GID>548</GID>
<name>OUT</name></connection>
<connection>
<GID>544</GID>
<name>IN_B_3</name></connection></vsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265.5,-63.5,265.5,-59.5</points>
<connection>
<GID>556</GID>
<name>IN_1</name></connection>
<connection>
<GID>552</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272,-63.5,272,-59.5</points>
<connection>
<GID>555</GID>
<name>IN_1</name></connection>
<connection>
<GID>551</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-63.5,277,-60</points>
<connection>
<GID>554</GID>
<name>IN_1</name></connection>
<connection>
<GID>550</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>283.5,-63.5,283.5,-60.5</points>
<connection>
<GID>553</GID>
<name>IN_1</name></connection>
<connection>
<GID>549</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307.5,-62.5,307.5,-43.5</points>
<connection>
<GID>545</GID>
<name>IN_1</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286,-43.5,309,-43.5</points>
<connection>
<GID>557</GID>
<name>OUT_0</name></connection>
<connection>
<GID>586</GID>
<name>IN_0</name></connection>
<intersection>307.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301,-62.5,301,-42.5</points>
<connection>
<GID>546</GID>
<name>IN_1</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286,-42.5,309,-42.5</points>
<connection>
<GID>557</GID>
<name>OUT_1</name></connection>
<connection>
<GID>586</GID>
<name>IN_1</name></connection>
<intersection>301 0</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,-62.5,295.5,-41.5</points>
<connection>
<GID>547</GID>
<name>IN_1</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286,-41.5,309,-41.5</points>
<connection>
<GID>557</GID>
<name>OUT_2</name></connection>
<connection>
<GID>586</GID>
<name>IN_2</name></connection>
<intersection>295.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,-62.5,288.5,-40.5</points>
<connection>
<GID>548</GID>
<name>IN_1</name></connection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286,-40.5,309,-40.5</points>
<connection>
<GID>557</GID>
<name>OUT_3</name></connection>
<connection>
<GID>586</GID>
<name>IN_3</name></connection>
<intersection>288.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-72,284.5,-69.5</points>
<connection>
<GID>558</GID>
<name>IN_1</name></connection>
<connection>
<GID>553</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-83,285.5,-78</points>
<connection>
<GID>558</GID>
<name>OUT</name></connection>
<connection>
<GID>544</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-72.5,278,-69.5</points>
<connection>
<GID>559</GID>
<name>IN_1</name></connection>
<connection>
<GID>554</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-83,284.5,-79.5</points>
<connection>
<GID>544</GID>
<name>IN_1</name></connection>
<intersection>-79.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>279,-79.5,284.5,-79.5</points>
<intersection>279 3</intersection>
<intersection>284.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>279,-79.5,279,-78.5</points>
<connection>
<GID>559</GID>
<name>OUT</name></connection>
<intersection>-79.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>283.5,-83,283.5,-80.5</points>
<connection>
<GID>544</GID>
<name>IN_2</name></connection>
<intersection>-80.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>274,-80.5,274,-78.5</points>
<connection>
<GID>560</GID>
<name>OUT</name></connection>
<intersection>-80.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>274,-80.5,283.5,-80.5</points>
<intersection>274 1</intersection>
<intersection>283.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282.5,-83,282.5,-81.5</points>
<connection>
<GID>544</GID>
<name>IN_3</name></connection>
<intersection>-81.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>267.5,-81.5,267.5,-78.5</points>
<connection>
<GID>561</GID>
<name>OUT</name></connection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>267.5,-81.5,282.5,-81.5</points>
<intersection>267.5 1</intersection>
<intersection>282.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273,-72.5,273,-69.5</points>
<connection>
<GID>560</GID>
<name>IN_1</name></connection>
<connection>
<GID>555</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266.5,-72.5,266.5,-69.5</points>
<connection>
<GID>561</GID>
<name>IN_1</name></connection>
<connection>
<GID>556</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268.5,-72.5,268.5,-71</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>265,-71,286.5,-71</points>
<connection>
<GID>562</GID>
<name>OUT_0</name></connection>
<intersection>268.5 0</intersection>
<intersection>275 3</intersection>
<intersection>280 5</intersection>
<intersection>286.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>275,-72.5,275,-71</points>
<connection>
<GID>560</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>280,-72.5,280,-71</points>
<connection>
<GID>559</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>286.5,-72,286.5,-71</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267.5,-63.5,267.5,-52.5</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,-52.5,316.5,-52.5</points>
<intersection>267.5 0</intersection>
<intersection>274 7</intersection>
<intersection>279 6</intersection>
<intersection>285.5 5</intersection>
<intersection>316.5 9</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>285.5,-63.5,285.5,-52.5</points>
<connection>
<GID>553</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>279,-63.5,279,-52.5</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>274,-63.5,274,-52.5</points>
<connection>
<GID>555</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>316.5,-62,316.5,-52.5</points>
<connection>
<GID>564</GID>
<name>IN_1</name></connection>
<intersection>-54.5 10</intersection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>316.5,-54.5,322.5,-54.5</points>
<connection>
<GID>597</GID>
<name>IN_0</name></connection>
<intersection>316.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-62.5,290.5,-51.5</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,-51.5,318.5,-51.5</points>
<intersection>290.5 0</intersection>
<intersection>297.5 3</intersection>
<intersection>303 7</intersection>
<intersection>309.5 6</intersection>
<intersection>318.5 9</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>297.5,-62.5,297.5,-51.5</points>
<connection>
<GID>547</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>309.5,-62.5,309.5,-51.5</points>
<connection>
<GID>545</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>303,-62.5,303,-51.5</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>318.5,-62,318.5,-51.5</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<intersection>-59 10</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>318.5,-59,324,-59</points>
<connection>
<GID>596</GID>
<name>IN_0</name></connection>
<intersection>318.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,-95.5,289,-91</points>
<connection>
<GID>544</GID>
<name>OUT_0</name></connection>
<intersection>-95.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>238,-95.5,289,-95.5</points>
<connection>
<GID>569</GID>
<name>IN_0</name></connection>
<intersection>246 8</intersection>
<intersection>289 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>246,-95.5,246,-85</points>
<connection>
<GID>573</GID>
<name>IN_3</name></connection>
<intersection>-95.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,-94,288,-91</points>
<connection>
<GID>544</GID>
<name>OUT_1</name></connection>
<intersection>-94 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>232.5,-94,288,-94</points>
<connection>
<GID>570</GID>
<name>IN_0</name></connection>
<intersection>244 8</intersection>
<intersection>288 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>244,-94,244,-85</points>
<connection>
<GID>573</GID>
<name>IN_2</name></connection>
<intersection>-94 7</intersection></vsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287,-92.5,287,-91</points>
<connection>
<GID>544</GID>
<name>OUT_2</name></connection>
<intersection>-92.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>239,-92.5,287,-92.5</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>242 8</intersection>
<intersection>287 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>242,-92.5,242,-85</points>
<connection>
<GID>573</GID>
<name>IN_1</name></connection>
<intersection>-92.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>233,-91,286,-91</points>
<connection>
<GID>544</GID>
<name>OUT_3</name></connection>
<connection>
<GID>572</GID>
<name>IN_0</name></connection>
<intersection>240 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>240,-91,240,-85</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>-91 7</intersection></vsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317.5,-86,317.5,-68</points>
<connection>
<GID>564</GID>
<name>OUT</name></connection>
<intersection>-86 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-86,317.5,-86</points>
<connection>
<GID>544</GID>
<name>carry_in</name></connection>
<intersection>317.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>273,-40.5,278,-40.5</points>
<connection>
<GID>531</GID>
<name>OUT_3</name></connection>
<connection>
<GID>557</GID>
<name>IN_3</name></connection>
<intersection>273 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>273,-40.5,273,-34.5</points>
<connection>
<GID>532</GID>
<name>OUT_0</name></connection>
<intersection>-40.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>273,-41.5,278,-41.5</points>
<connection>
<GID>531</GID>
<name>OUT_2</name></connection>
<connection>
<GID>557</GID>
<name>IN_2</name></connection>
<intersection>274 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>274,-41.5,274,-34.5</points>
<connection>
<GID>532</GID>
<name>OUT_1</name></connection>
<intersection>-41.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>273,-42.5,278,-42.5</points>
<connection>
<GID>531</GID>
<name>OUT_1</name></connection>
<connection>
<GID>557</GID>
<name>IN_1</name></connection>
<intersection>275 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>275,-42.5,275,-34.5</points>
<connection>
<GID>532</GID>
<name>OUT_2</name></connection>
<intersection>-42.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>273,-43.5,278,-43.5</points>
<connection>
<GID>531</GID>
<name>OUT_0</name></connection>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<intersection>276 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>276,-43.5,276,-34.5</points>
<connection>
<GID>532</GID>
<name>OUT_3</name></connection>
<intersection>-43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,-40.5,269,-40.5</points>
<connection>
<GID>531</GID>
<name>IN_3</name></connection>
<connection>
<GID>533</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>261.5,-41.5,269,-41.5</points>
<connection>
<GID>531</GID>
<name>IN_2</name></connection>
<connection>
<GID>534</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>256,-42.5,269,-42.5</points>
<connection>
<GID>531</GID>
<name>IN_1</name></connection>
<connection>
<GID>535</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>250,-43.5,269,-43.5</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<connection>
<GID>536</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-30.5,276,-29.5</points>
<connection>
<GID>532</GID>
<name>IN_3</name></connection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>276,-29.5,323.5,-29.5</points>
<intersection>276 0</intersection>
<intersection>318.5 4</intersection>
<intersection>323.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>323.5,-29.5,323.5,-25.5</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<intersection>-29.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>318.5,-43.5,318.5,-29.5</points>
<intersection>-43.5 5</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>313,-43.5,318.5,-43.5</points>
<connection>
<GID>586</GID>
<name>OUT_0</name></connection>
<intersection>318.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319.5,-28.5,319.5,-25</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<intersection>-28.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>275,-28.5,319.5,-28.5</points>
<intersection>275 8</intersection>
<intersection>316 9</intersection>
<intersection>319.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>275,-30.5,275,-28.5</points>
<connection>
<GID>532</GID>
<name>IN_2</name></connection>
<intersection>-28.5 7</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>316,-42.5,316,-28.5</points>
<intersection>-42.5 10</intersection>
<intersection>-28.5 7</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>313,-42.5,316,-42.5</points>
<connection>
<GID>586</GID>
<name>OUT_1</name></connection>
<intersection>316 9</intersection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-30.5,274,-27.5</points>
<connection>
<GID>532</GID>
<name>IN_1</name></connection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>274,-27.5,316.5,-27.5</points>
<intersection>274 0</intersection>
<intersection>314.5 8</intersection>
<intersection>316.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>316.5,-27.5,316.5,-25</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<intersection>-27.5 3</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>314.5,-41.5,314.5,-27.5</points>
<intersection>-41.5 9</intersection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>313,-41.5,314.5,-41.5</points>
<connection>
<GID>586</GID>
<name>OUT_2</name></connection>
<intersection>314.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273,-30.5,273,-26</points>
<connection>
<GID>532</GID>
<name>IN_0</name></connection>
<intersection>-26 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>313,-40.5,313,-24.5</points>
<connection>
<GID>586</GID>
<name>OUT_3</name></connection>
<connection>
<GID>540</GID>
<name>IN_0</name></connection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>273,-26,313,-26</points>
<intersection>273 0</intersection>
<intersection>313 1</intersection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-48,281,-46.5</points>
<connection>
<GID>557</GID>
<name>clock</name></connection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277.5,-48,281,-48</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>283,-46.5,283,-46.5</points>
<connection>
<GID>542</GID>
<name>OUT_0</name></connection>
<connection>
<GID>557</GID>
<name>clear</name></connection></hsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-37.5,282,-36</points>
<connection>
<GID>557</GID>
<name>count_enable</name></connection>
<connection>
<GID>543</GID>
<name>OUT_0</name></connection>
<intersection>-37 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>282,-37,283,-37</points>
<intersection>282 0</intersection>
<intersection>283 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>283,-37.5,283,-37</points>
<connection>
<GID>557</GID>
<name>count_up</name></connection>
<intersection>-37 3</intersection></vsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-37.5,281,-33</points>
<connection>
<GID>557</GID>
<name>load</name></connection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281,-33,290,-33</points>
<connection>
<GID>567</GID>
<name>IN_0</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>256,-71,261,-71</points>
<connection>
<GID>562</GID>
<name>IN_0</name></connection>
<connection>
<GID>568</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-78,243,-73</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<connection>
<GID>573</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118,-86,191.5,-86</points>
<connection>
<GID>431</GID>
<name>carry_in</name></connection>
<connection>
<GID>498</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>207.5,-86,279.5,-86</points>
<connection>
<GID>498</GID>
<name>carry_in</name></connection>
<connection>
<GID>544</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-39,311,-38</points>
<connection>
<GID>586</GID>
<name>ENABLE_0</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309,-38,311,-38</points>
<connection>
<GID>588</GID>
<name>IN_0</name></connection>
<intersection>311 0</intersection></hsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,-39,222.5,-37.5</points>
<connection>
<GID>589</GID>
<name>ENABLE_0</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>220.5,-37.5,222.5,-37.5</points>
<connection>
<GID>590</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,-39,133.5,-37.5</points>
<connection>
<GID>591</GID>
<name>ENABLE_0</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-37.5,133.5,-37.5</points>
<connection>
<GID>592</GID>
<name>IN_0</name></connection>
<intersection>133.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-40,42,-38.5</points>
<connection>
<GID>593</GID>
<name>ENABLE_0</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-38.5,42,-38.5</points>
<connection>
<GID>594</GID>
<name>IN_0</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-38.5,13,-37</points>
<connection>
<GID>369</GID>
<name>load</name></connection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-37,13,-37</points>
<connection>
<GID>608</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59.5,-34,-59.5,-29.5</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<connection>
<GID>519</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,-34,-56.5,-32</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-57.5,-32,-57.5,-29.5</points>
<connection>
<GID>519</GID>
<name>IN_1</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,-32,-56.5,-32</points>
<intersection>-57.5 1</intersection>
<intersection>-56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-34.5,-52,-32</points>
<connection>
<GID>603</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-55.5,-32,-55.5,-29.5</points>
<connection>
<GID>519</GID>
<name>IN_2</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-55.5,-32,-52,-32</points>
<intersection>-55.5 1</intersection>
<intersection>-52 0</intersection></hsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-34.5,-49,-31</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-53.5,-31,-53.5,-29.5</points>
<connection>
<GID>519</GID>
<name>IN_3</name></connection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-53.5,-31,-49,-31</points>
<intersection>-53.5 1</intersection>
<intersection>-49 0</intersection></hsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,-17.5,-56.5,-16</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<connection>
<GID>529</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>630</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,-23.5,-56.5,-22.5</points>
<connection>
<GID>519</GID>
<name>OUT</name></connection>
<intersection>-22.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-57.5,-22.5,-57.5,-21.5</points>
<connection>
<GID>529</GID>
<name>IN_1</name></connection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,-22.5,-56.5,-22.5</points>
<intersection>-57.5 1</intersection>
<intersection>-56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>631</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-63,-19.5,-59,-19.5</points>
<connection>
<GID>529</GID>
<name>SEL_0</name></connection>
<connection>
<GID>563</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>632</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-65,-68.5,-61,-68.5</points>
<connection>
<GID>565</GID>
<name>SEL_0</name></connection>
<connection>
<GID>566</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>661</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-96.5,21,-92</points>
<connection>
<GID>335</GID>
<name>OUT_0</name></connection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63,-96.5,21,-96.5</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>-34.5 2</intersection>
<intersection>21 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-34.5,-96.5,-34.5,-86.5</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>-96.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>662</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54,-64,-54,-62</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>-64 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-58.5,-66.5,-58.5,-64</points>
<connection>
<GID>565</GID>
<name>OUT</name></connection>
<intersection>-64 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-58.5,-64,-54,-64</points>
<intersection>-58.5 1</intersection>
<intersection>-54 0</intersection></hsegment></shape></wire>
<wire>
<ID>668</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-83.5,-46.5,-83.5</points>
<connection>
<GID>575</GID>
<name>SEL_0</name></connection>
<connection>
<GID>576</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>669</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-81.5,-44,-81</points>
<connection>
<GID>575</GID>
<name>OUT</name></connection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-44,-81,-43,-81</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-84,40.5,-69.5</points>
<connection>
<GID>338</GID>
<name>OUT</name></connection>
<intersection>-84 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-84,40.5,-84</points>
<connection>
<GID>335</GID>
<name>IN_B_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-83,34,-69.5</points>
<connection>
<GID>339</GID>
<name>OUT</name></connection>
<intersection>-83 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>23.5,-83,34,-83</points>
<intersection>23.5 4</intersection>
<intersection>34 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>23.5,-84,23.5,-83</points>
<connection>
<GID>335</GID>
<name>IN_B_1</name></connection>
<intersection>-83 3</intersection></vsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-84,22.5,-82</points>
<connection>
<GID>335</GID>
<name>IN_B_2</name></connection>
<intersection>-82 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>28.5,-82,28.5,-69.5</points>
<connection>
<GID>340</GID>
<name>OUT</name></connection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-82,28.5,-82</points>
<intersection>22.5 0</intersection>
<intersection>28.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-84,21.5,-69.5</points>
<connection>
<GID>341</GID>
<name>OUT</name></connection>
<connection>
<GID>335</GID>
<name>IN_B_3</name></connection></vsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,-78,-45,-78</points>
<connection>
<GID>337</GID>
<name>OUT_0</name></connection>
<connection>
<GID>336</GID>
<name>set</name></connection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-37,-78,-32,-78</points>
<connection>
<GID>336</GID>
<name>clear</name></connection>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>-40,-81.5,-40,-81</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<connection>
<GID>336</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-86.5,-36.5,-73.5</points>
<intersection>-86.5 8</intersection>
<intersection>-73.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-44,-73.5,-36.5,-73.5</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>-43 11</intersection>
<intersection>-36.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-43,-86.5,-36.5,-86.5</points>
<intersection>-43 12</intersection>
<intersection>-36.5 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-43,-75,-43,-71.5</points>
<connection>
<GID>336</GID>
<name>OUT_0</name></connection>
<connection>
<GID>349</GID>
<name>N_in2</name></connection>
<intersection>-73.5 6</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-43,-86.5,-43,-85.5</points>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<intersection>-86.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-25.5,-77.5,-24.5,-77.5</points>
<connection>
<GID>356</GID>
<name>set</name></connection>
<connection>
<GID>357</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16.5,-77.5,-14,-77.5</points>
<connection>
<GID>356</GID>
<name>clear</name></connection>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>-19.5,-81,-19.5,-80.5</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<connection>
<GID>356</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-86,-11,-72.5</points>
<intersection>-86 14</intersection>
<intersection>-72.5 15</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-21.5,-86,-11,-86</points>
<intersection>-21.5 19</intersection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-22.5,-72.5,-11,-72.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>-22.5 18</intersection>
<intersection>-11 0</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>-22.5,-74.5,-22.5,-71</points>
<connection>
<GID>360</GID>
<name>N_in2</name></connection>
<connection>
<GID>356</GID>
<name>OUT_0</name></connection>
<intersection>-72.5 15</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>-21.5,-86,-21.5,-84.5</points>
<connection>
<GID>577</GID>
<name>IN_0</name></connection>
<intersection>-86 14</intersection></vsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-57,-59,-56,-59</points>
<connection>
<GID>366</GID>
<name>OUT_0</name></connection>
<connection>
<GID>364</GID>
<name>set</name></connection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48,-59,-47,-59</points>
<connection>
<GID>368</GID>
<name>OUT_0</name></connection>
<connection>
<GID>364</GID>
<name>clear</name></connection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>14</ID>
<points>-51,-62.5,-51,-62</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<connection>
<GID>364</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>692</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45,-87,-45,-85.5</points>
<connection>
<GID>575</GID>
<name>IN_1</name></connection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49,-87,11.5,-87</points>
<connection>
<GID>335</GID>
<name>carry_out</name></connection>
<connection>
<GID>350</GID>
<name>N_in1</name></connection>
<intersection>-45 0</intersection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,-70.5,-44.5,-54.5</points>
<intersection>-70.5 7</intersection>
<intersection>-54.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-55,-54.5,-44.5,-54.5</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>-54 10</intersection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-57.5,-70.5,-44.5,-70.5</points>
<connection>
<GID>565</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-54,-56,-54,-52.5</points>
<connection>
<GID>364</GID>
<name>OUT_0</name></connection>
<connection>
<GID>375</GID>
<name>N_in2</name></connection>
<intersection>-54.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-58.5,-13,-57.5,-13</points>
<connection>
<GID>379</GID>
<name>set</name></connection>
<intersection>-57.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-57.5,-13,-57.5,-12</points>
<connection>
<GID>381</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-50.5,-13,-47.5,-13</points>
<connection>
<GID>379</GID>
<name>clear</name></connection>
<intersection>-47.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-47.5,-13,-47.5,-12</points>
<connection>
<GID>383</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-64.5,-2.5,-60.5</points>
<connection>
<GID>354</GID>
<name>IN_1</name></connection>
<connection>
<GID>346</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-64.5,4,-62.5</points>
<connection>
<GID>353</GID>
<name>IN_1</name></connection>
<connection>
<GID>345</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-64.5,9,-62</points>
<connection>
<GID>352</GID>
<name>IN_1</name></connection>
<connection>
<GID>344</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-64.5,15.5,-63</points>
<connection>
<GID>351</GID>
<name>IN_1</name></connection>
<connection>
<GID>343</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>12</ID>
<points>-52,-17.5,-52,-16</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>-16 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-53.5,-16,-52,-16</points>
<connection>
<GID>379</GID>
<name>clock</name></connection>
<intersection>-52 12</intersection></hsegment></shape></wire>
<wire>
<ID>702</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>-25,-82.5,-25,-68.5</points>
<connection>
<GID>577</GID>
<name>SEL_0</name></connection>
<intersection>-68.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-30.5,-68.5,-25,-68.5</points>
<connection>
<GID>578</GID>
<name>IN_0</name></connection>
<intersection>-25 4</intersection></hsegment></shape></wire>
<wire>
<ID>703</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-80.5,-22.5,-80.5</points>
<connection>
<GID>577</GID>
<name>OUT</name></connection>
<connection>
<GID>356</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>704</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23.5,-89,-23.5,-84.5</points>
<connection>
<GID>577</GID>
<name>IN_1</name></connection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-89,11.5,-89</points>
<connection>
<GID>335</GID>
<name>overflow</name></connection>
<connection>
<GID>347</GID>
<name>N_in1</name></connection>
<intersection>-23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43.5,-23,-43.5,-7.5</points>
<intersection>-23 7</intersection>
<intersection>-7.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-58,-7.5,-43.5,-7.5</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>-56.5 11</intersection>
<intersection>-43.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-55.5,-23,-43.5,-23</points>
<intersection>-55.5 10</intersection>
<intersection>-43.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-55.5,-23,-55.5,-21.5</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>-23 7</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-56.5,-10,-56.5,-5.5</points>
<connection>
<GID>379</GID>
<name>OUT_0</name></connection>
<connection>
<GID>389</GID>
<name>N_in2</name></connection>
<intersection>-7.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-63.5,39.5,-44.5</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-44.5,40,-44.5</points>
<connection>
<GID>369</GID>
<name>OUT_0</name></connection>
<connection>
<GID>593</GID>
<name>IN_0</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-63.5,33,-43.5</points>
<connection>
<GID>339</GID>
<name>IN_1</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-43.5,40,-43.5</points>
<connection>
<GID>369</GID>
<name>OUT_1</name></connection>
<connection>
<GID>593</GID>
<name>IN_1</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-63.5,27.5,-42.5</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-42.5,40,-42.5</points>
<connection>
<GID>369</GID>
<name>OUT_2</name></connection>
<connection>
<GID>593</GID>
<name>IN_2</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-63.5,20.5,-41.5</points>
<connection>
<GID>341</GID>
<name>IN_1</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-41.5,40,-41.5</points>
<connection>
<GID>369</GID>
<name>OUT_3</name></connection>
<connection>
<GID>593</GID>
<name>IN_3</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-73,16.5,-70.5</points>
<connection>
<GID>371</GID>
<name>IN_1</name></connection>
<connection>
<GID>351</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-84,17.5,-79</points>
<connection>
<GID>371</GID>
<name>OUT</name></connection>
<connection>
<GID>335</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-73.5,10,-70.5</points>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<connection>
<GID>352</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-84,16.5,-80.5</points>
<connection>
<GID>335</GID>
<name>IN_1</name></connection>
<intersection>-80.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>11,-80.5,11,-79.5</points>
<connection>
<GID>372</GID>
<name>OUT</name></connection>
<intersection>-80.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11,-80.5,16.5,-80.5</points>
<intersection>11 1</intersection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-84,15.5,-81.5</points>
<connection>
<GID>335</GID>
<name>IN_2</name></connection>
<intersection>-81.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>6,-81.5,6,-79.5</points>
<connection>
<GID>373</GID>
<name>OUT</name></connection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>6,-81.5,15.5,-81.5</points>
<intersection>6 1</intersection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-84,14.5,-82.5</points>
<connection>
<GID>335</GID>
<name>IN_3</name></connection>
<intersection>-82.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-0.5,-82.5,-0.5,-79.5</points>
<connection>
<GID>374</GID>
<name>OUT</name></connection>
<intersection>-82.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,-82.5,14.5,-82.5</points>
<intersection>-0.5 1</intersection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-73.5,5,-70.5</points>
<connection>
<GID>373</GID>
<name>IN_1</name></connection>
<connection>
<GID>353</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-73.5,-1.5,-70.5</points>
<connection>
<GID>374</GID>
<name>IN_1</name></connection>
<connection>
<GID>354</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-73.5,0.5,-72</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3,-72,18.5,-72</points>
<connection>
<GID>376</GID>
<name>OUT_0</name></connection>
<intersection>0.5 0</intersection>
<intersection>7 3</intersection>
<intersection>12 5</intersection>
<intersection>18.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>7,-73.5,7,-72</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>-72 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>12,-73.5,12,-72</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>-72 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>18.5,-73,18.5,-72</points>
<connection>
<GID>371</GID>
<name>IN_0</name></connection>
<intersection>-72 1</intersection></vsegment></shape></wire>
<wire>
<ID>719</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,-6,289,-4.86719e-008</points>
<connection>
<GID>660</GID>
<name>OUT_0</name></connection>
<connection>
<GID>479</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-64.5,-0.5,-51.5</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-51.5,47,-51.5</points>
<connection>
<GID>606</GID>
<name>IN_0</name></connection>
<intersection>-0.5 0</intersection>
<intersection>6 7</intersection>
<intersection>11 6</intersection>
<intersection>17.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>17.5,-64.5,17.5,-51.5</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>11,-64.5,11,-51.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>6,-64.5,6,-51.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-63.5,22.5,-52.5</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-52.5,41.5,-52.5</points>
<intersection>22.5 0</intersection>
<intersection>29.5 3</intersection>
<intersection>35 7</intersection>
<intersection>41.5 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>29.5,-63.5,29.5,-52.5</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>41.5,-63.5,41.5,-52.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>-55.5 10</intersection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>35,-63.5,35,-52.5</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>41.5,-55.5,49,-55.5</points>
<connection>
<GID>605</GID>
<name>IN_0</name></connection>
<intersection>41.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-95,20,-92</points>
<connection>
<GID>335</GID>
<name>OUT_1</name></connection>
<intersection>-95 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-68.5,-95,20,-95</points>
<connection>
<GID>391</GID>
<name>IN_0</name></connection>
<intersection>-32.5 13</intersection>
<intersection>20 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-32.5,-95,-32.5,-86.5</points>
<connection>
<GID>397</GID>
<name>IN_1</name></connection>
<intersection>-95 8</intersection></vsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-93.5,19,-92</points>
<connection>
<GID>335</GID>
<name>OUT_2</name></connection>
<intersection>-93.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-62,-93.5,19,-93.5</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>-30.5 13</intersection>
<intersection>19 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-30.5,-93.5,-30.5,-86.5</points>
<connection>
<GID>397</GID>
<name>IN_2</name></connection>
<intersection>-93.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-68,-92,18,-92</points>
<connection>
<GID>335</GID>
<name>OUT_3</name></connection>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<intersection>-59.5 16</intersection>
<intersection>-28.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-28.5,-92,-28.5,-86.5</points>
<connection>
<GID>397</GID>
<name>IN_3</name></connection>
<intersection>-92 10</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-59.5,-92,-59.5,-70.5</points>
<connection>
<GID>565</GID>
<name>IN_1</name></connection>
<intersection>-92 10</intersection></vsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-41.5,10,-41.5</points>
<connection>
<GID>369</GID>
<name>IN_3</name></connection>
<connection>
<GID>395</GID>
<name>OUT_3</name></connection>
<intersection>5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>5,-41.5,5,-35.5</points>
<connection>
<GID>396</GID>
<name>OUT_0</name></connection>
<intersection>-41.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-42.5,10,-42.5</points>
<connection>
<GID>369</GID>
<name>IN_2</name></connection>
<connection>
<GID>395</GID>
<name>OUT_2</name></connection>
<intersection>6 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>6,-42.5,6,-35.5</points>
<connection>
<GID>396</GID>
<name>OUT_1</name></connection>
<intersection>-42.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-43.5,10,-43.5</points>
<connection>
<GID>369</GID>
<name>IN_1</name></connection>
<connection>
<GID>395</GID>
<name>OUT_1</name></connection>
<intersection>7 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>7,-43.5,7,-35.5</points>
<connection>
<GID>396</GID>
<name>OUT_2</name></connection>
<intersection>-43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5,-44.5,10,-44.5</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<connection>
<GID>395</GID>
<name>OUT_0</name></connection>
<intersection>8 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>8,-44.5,8,-35.5</points>
<connection>
<GID>396</GID>
<name>OUT_3</name></connection>
<intersection>-44.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-41.5,1,-41.5</points>
<connection>
<GID>395</GID>
<name>IN_3</name></connection>
<connection>
<GID>398</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-6.5,-42.5,1,-42.5</points>
<connection>
<GID>395</GID>
<name>IN_2</name></connection>
<connection>
<GID>399</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-43.5,1,-43.5</points>
<connection>
<GID>395</GID>
<name>IN_1</name></connection>
<connection>
<GID>400</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18,-44.5,1,-44.5</points>
<connection>
<GID>395</GID>
<name>IN_0</name></connection>
<connection>
<GID>401</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-31.5,8,-30</points>
<connection>
<GID>396</GID>
<name>IN_3</name></connection>
<intersection>-30 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>55,-44.5,55,-24.5</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<intersection>-44.5 4</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>8,-30,55,-30</points>
<intersection>8 0</intersection>
<intersection>55 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>44,-44.5,55,-44.5</points>
<connection>
<GID>593</GID>
<name>OUT_0</name></connection>
<intersection>55 1</intersection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-43.5,51,-24</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<intersection>-43.5 6</intersection>
<intersection>-28.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>7,-28.5,51,-28.5</points>
<intersection>7 4</intersection>
<intersection>51 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>7,-31.5,7,-28.5</points>
<connection>
<GID>396</GID>
<name>IN_2</name></connection>
<intersection>-28.5 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>44,-43.5,51,-43.5</points>
<connection>
<GID>593</GID>
<name>OUT_1</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-31.5,6,-27.5</points>
<connection>
<GID>396</GID>
<name>IN_1</name></connection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>6,-27.5,47,-27.5</points>
<intersection>6 0</intersection>
<intersection>47 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>47,-42.5,47,-23.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<intersection>-42.5 7</intersection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>44,-42.5,47,-42.5</points>
<connection>
<GID>593</GID>
<name>OUT_2</name></connection>
<intersection>47 5</intersection></hsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-31.5,5,-25.5</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>44,-41.5,44,-23.5</points>
<connection>
<GID>593</GID>
<name>OUT_3</name></connection>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>5,-25.5,44,-25.5</points>
<intersection>5 0</intersection>
<intersection>44 1</intersection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-49,13,-47.5</points>
<connection>
<GID>369</GID>
<name>clock</name></connection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,-49,13,-49</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-47.5,15,-47.5</points>
<connection>
<GID>407</GID>
<name>OUT_0</name></connection>
<connection>
<GID>369</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-38.5,14,-36.5</points>
<connection>
<GID>369</GID>
<name>count_enable</name></connection>
<connection>
<GID>408</GID>
<name>OUT_0</name></connection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>14,-38.5,15,-38.5</points>
<connection>
<GID>369</GID>
<name>count_up</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-83,131,-68.5</points>
<connection>
<GID>432</GID>
<name>OUT</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-83,131,-83</points>
<connection>
<GID>431</GID>
<name>IN_B_0</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-82,124.5,-68.5</points>
<connection>
<GID>433</GID>
<name>OUT</name></connection>
<intersection>-82 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>114,-82,124.5,-82</points>
<intersection>114 4</intersection>
<intersection>124.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>114,-83,114,-82</points>
<connection>
<GID>431</GID>
<name>IN_B_1</name></connection>
<intersection>-82 3</intersection></vsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-83,113,-81</points>
<connection>
<GID>431</GID>
<name>IN_B_2</name></connection>
<intersection>-81 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>119,-81,119,-68.5</points>
<connection>
<GID>434</GID>
<name>OUT</name></connection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>113,-81,119,-81</points>
<intersection>113 0</intersection>
<intersection>119 1</intersection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-83,112,-68.5</points>
<connection>
<GID>431</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>435</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9.5,-33.5,16,-33.5</points>
<connection>
<GID>396</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>382</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-32.5,100,-32.5</points>
<connection>
<GID>419</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>384</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-63.5,88,-59.5</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<connection>
<GID>443</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,-63.5,94.5,-59.5</points>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<connection>
<GID>442</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-63.5,99.5,-60</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<connection>
<GID>441</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-63.5,106,-60.5</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<connection>
<GID>440</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-62.5,130,-43.5</points>
<connection>
<GID>432</GID>
<name>IN_1</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-43.5,131.5,-43.5</points>
<connection>
<GID>450</GID>
<name>OUT_0</name></connection>
<connection>
<GID>591</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-62.5,123.5,-42.5</points>
<connection>
<GID>433</GID>
<name>IN_1</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-42.5,131.5,-42.5</points>
<connection>
<GID>450</GID>
<name>OUT_1</name></connection>
<connection>
<GID>591</GID>
<name>IN_1</name></connection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-62.5,118,-41.5</points>
<connection>
<GID>434</GID>
<name>IN_1</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-41.5,131.5,-41.5</points>
<connection>
<GID>450</GID>
<name>OUT_2</name></connection>
<connection>
<GID>591</GID>
<name>IN_2</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-62.5,111,-40.5</points>
<connection>
<GID>435</GID>
<name>IN_1</name></connection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-40.5,131.5,-40.5</points>
<connection>
<GID>450</GID>
<name>OUT_3</name></connection>
<connection>
<GID>591</GID>
<name>IN_3</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-72,107,-69.5</points>
<connection>
<GID>440</GID>
<name>OUT</name></connection>
<connection>
<GID>451</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-83,108,-78</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<connection>
<GID>451</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-72.5,100.5,-69.5</points>
<connection>
<GID>441</GID>
<name>OUT</name></connection>
<connection>
<GID>452</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-83,107,-79.5</points>
<connection>
<GID>431</GID>
<name>IN_1</name></connection>
<intersection>-79.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>101.5,-79.5,107,-79.5</points>
<intersection>101.5 3</intersection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>101.5,-79.5,101.5,-78.5</points>
<connection>
<GID>452</GID>
<name>OUT</name></connection>
<intersection>-79.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-83,106,-80.5</points>
<connection>
<GID>431</GID>
<name>IN_2</name></connection>
<intersection>-80.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>96.5,-80.5,96.5,-78.5</points>
<connection>
<GID>453</GID>
<name>OUT</name></connection>
<intersection>-80.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-80.5,106,-80.5</points>
<intersection>96.5 1</intersection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-83,105,-81.5</points>
<connection>
<GID>431</GID>
<name>IN_3</name></connection>
<intersection>-81.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>90,-81.5,90,-78.5</points>
<connection>
<GID>454</GID>
<name>OUT</name></connection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>90,-81.5,105,-81.5</points>
<intersection>90 1</intersection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-72.5,95.5,-69.5</points>
<connection>
<GID>442</GID>
<name>OUT</name></connection>
<connection>
<GID>453</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-72.5,89,-69.5</points>
<connection>
<GID>443</GID>
<name>OUT</name></connection>
<connection>
<GID>454</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-72.5,91,-71</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87.5,-71,109,-71</points>
<connection>
<GID>455</GID>
<name>OUT_0</name></connection>
<intersection>91 0</intersection>
<intersection>97.5 3</intersection>
<intersection>102.5 5</intersection>
<intersection>109 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>97.5,-72.5,97.5,-71</points>
<connection>
<GID>453</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>102.5,-72.5,102.5,-71</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>109,-72,109,-71</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<intersection>-71 1</intersection></vsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-63.5,90,-52.5</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-52.5,108,-52.5</points>
<intersection>90 0</intersection>
<intersection>96.5 7</intersection>
<intersection>101.5 6</intersection>
<intersection>108 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>108,-63.5,108,-52.5</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<intersection>-53.5 10</intersection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>101.5,-63.5,101.5,-52.5</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>96.5,-63.5,96.5,-52.5</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>108,-53.5,136,-53.5</points>
<connection>
<GID>602</GID>
<name>IN_0</name></connection>
<intersection>108 5</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-249.478,178.648,876.522,-467.352</PageViewport>
<gate>
<ID>3</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-65,-5</position>
<input>
<ID>ENABLE_0</ID>179 </input>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>84 </input>
<input>
<ID>IN_2</ID>83 </input>
<input>
<ID>IN_3</ID>82 </input>
<input>
<ID>IN_4</ID>81 </input>
<input>
<ID>IN_5</ID>80 </input>
<input>
<ID>IN_6</ID>79 </input>
<input>
<ID>IN_7</ID>78 </input>
<output>
<ID>OUT_0</ID>178 </output>
<output>
<ID>OUT_1</ID>177 </output>
<output>
<ID>OUT_2</ID>176 </output>
<output>
<ID>OUT_3</ID>130 </output>
<output>
<ID>OUT_4</ID>93 </output>
<output>
<ID>OUT_5</ID>92 </output>
<output>
<ID>OUT_6</ID>91 </output>
<output>
<ID>OUT_7</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>7</ID>
<type>DE_TO</type>
<position>-60.5,8.5</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I11</lparam></gate>
<gate>
<ID>9</ID>
<type>DE_TO</type>
<position>-60.5,6.5</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I10</lparam></gate>
<gate>
<ID>11</ID>
<type>DE_TO</type>
<position>-60.5,4</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I9</lparam></gate>
<gate>
<ID>13</ID>
<type>DE_TO</type>
<position>-60.5,2</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I8</lparam></gate>
<gate>
<ID>15</ID>
<type>DE_TO</type>
<position>-49.5,-1.5</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I7</lparam></gate>
<gate>
<ID>17</ID>
<type>DE_TO</type>
<position>-49.5,-3.5</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I6</lparam></gate>
<gate>
<ID>19</ID>
<type>DE_TO</type>
<position>-49.5,-6</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I5</lparam></gate>
<gate>
<ID>21</ID>
<type>DE_TO</type>
<position>-49.5,-8</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I4</lparam></gate>
<gate>
<ID>23</ID>
<type>DE_TO</type>
<position>-55.5,-10.5</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I3</lparam></gate>
<gate>
<ID>25</ID>
<type>DE_TO</type>
<position>-55.5,-12.5</position>
<input>
<ID>IN_0</ID>176 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I2</lparam></gate>
<gate>
<ID>803</ID>
<type>DA_FROM</type>
<position>-77,-1</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>804</ID>
<type>DA_FROM</type>
<position>-76.5,-3.5</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>805</ID>
<type>DA_FROM</type>
<position>-77.5,-6.5</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>806</ID>
<type>DA_FROM</type>
<position>-76.5,-9.5</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>807</ID>
<type>DA_FROM</type>
<position>-76.5,-11.5</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>808</ID>
<type>DA_FROM</type>
<position>-76.5,-14.5</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>809</ID>
<type>DA_FROM</type>
<position>-77,-17.5</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>-55.5,-15</position>
<input>
<ID>IN_0</ID>177 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I1</lparam></gate>
<gate>
<ID>810</ID>
<type>DA_FROM</type>
<position>-77,-21.5</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>812</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>-69,7</position>
<input>
<ID>ENABLE_0</ID>179 </input>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>45 </input>
<input>
<ID>IN_2</ID>4 </input>
<input>
<ID>IN_3</ID>701 </input>
<output>
<ID>OUT_0</ID>89 </output>
<output>
<ID>OUT_1</ID>88 </output>
<output>
<ID>OUT_2</ID>87 </output>
<output>
<ID>OUT_3</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>-55.5,-17</position>
<input>
<ID>IN_0</ID>178 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I0</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>-81.5,20.5</position>
<input>
<ID>IN_0</ID>179 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BUS-PC</lparam></gate>
<gate>
<ID>60</ID>
<type>DA_FROM</type>
<position>-15.5,-10.5</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I8</lparam></gate>
<gate>
<ID>61</ID>
<type>DA_FROM</type>
<position>-18,-10.5</position>
<input>
<ID>IN_0</ID>181 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I9</lparam></gate>
<gate>
<ID>62</ID>
<type>DA_FROM</type>
<position>-20.5,-10.5</position>
<input>
<ID>IN_0</ID>182 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I10</lparam></gate>
<gate>
<ID>65</ID>
<type>DA_FROM</type>
<position>-23,-10.5</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I11</lparam></gate>
<gate>
<ID>67</ID>
<type>DA_FROM</type>
<position>5,-11</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I4</lparam></gate>
<gate>
<ID>69</ID>
<type>DA_FROM</type>
<position>2.5,-11</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I5</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>0,-11</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I6</lparam></gate>
<gate>
<ID>74</ID>
<type>DA_FROM</type>
<position>-2.5,-11</position>
<input>
<ID>IN_0</ID>184 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I7</lparam></gate>
<gate>
<ID>275</ID>
<type>AA_TOGGLE</type>
<position>-9,-57.5</position>
<output>
<ID>OUT_0</ID>249 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>276</ID>
<type>DE_TO</type>
<position>-1,-57.5</position>
<input>
<ID>IN_0</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck3</lparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>25.5,-10.5</position>
<input>
<ID>IN_0</ID>192 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I0</lparam></gate>
<gate>
<ID>91</ID>
<type>DA_FROM</type>
<position>23,-10.5</position>
<input>
<ID>IN_0</ID>191 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I1</lparam></gate>
<gate>
<ID>675</ID>
<type>AA_LABEL</type>
<position>-46.5,33</position>
<gparam>LABEL_TEXT Program Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>677</ID>
<type>AI_REGISTER12</type>
<position>54.5,-39.5</position>
<input>
<ID>IN_0</ID>649 </input>
<input>
<ID>IN_1</ID>650 </input>
<input>
<ID>IN_10</ID>659 </input>
<input>
<ID>IN_11</ID>660 </input>
<input>
<ID>IN_2</ID>651 </input>
<input>
<ID>IN_3</ID>652 </input>
<input>
<ID>IN_4</ID>653 </input>
<input>
<ID>IN_5</ID>654 </input>
<input>
<ID>IN_6</ID>655 </input>
<input>
<ID>IN_7</ID>656 </input>
<input>
<ID>IN_8</ID>657 </input>
<input>
<ID>IN_9</ID>658 </input>
<output>
<ID>OUT_0</ID>603 </output>
<output>
<ID>OUT_1</ID>602 </output>
<output>
<ID>OUT_10</ID>596 </output>
<output>
<ID>OUT_11</ID>595 </output>
<output>
<ID>OUT_2</ID>601 </output>
<output>
<ID>OUT_3</ID>604 </output>
<output>
<ID>OUT_4</ID>600 </output>
<output>
<ID>OUT_5</ID>597 </output>
<output>
<ID>OUT_6</ID>594 </output>
<output>
<ID>OUT_7</ID>599 </output>
<output>
<ID>OUT_8</ID>598 </output>
<output>
<ID>OUT_9</ID>593 </output>
<input>
<ID>clear</ID>589 </input>
<input>
<ID>clock</ID>588 </input>
<input>
<ID>count_enable</ID>592 </input>
<input>
<ID>count_up</ID>590 </input>
<input>
<ID>load</ID>591 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>679</ID>
<type>DA_FROM</type>
<position>53.5,-51</position>
<input>
<ID>IN_0</ID>588 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>681</ID>
<type>DA_FROM</type>
<position>55.5,-53.5</position>
<input>
<ID>IN_0</ID>589 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>683</ID>
<type>EE_VDD</type>
<position>55.5,-28.5</position>
<output>
<ID>OUT_0</ID>590 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>685</ID>
<type>DA_FROM</type>
<position>48,-30</position>
<input>
<ID>IN_0</ID>591 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load PC</lparam></gate>
<gate>
<ID>687</ID>
<type>DA_FROM</type>
<position>47.5,-24.5</position>
<input>
<ID>IN_0</ID>592 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>109</ID>
<type>DA_FROM</type>
<position>20.5,-10.5</position>
<input>
<ID>IN_0</ID>190 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I2</lparam></gate>
<gate>
<ID>689</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>103,-37.5</position>
<input>
<ID>ENABLE_0</ID>605 </input>
<input>
<ID>IN_0</ID>600 </input>
<input>
<ID>IN_1</ID>597 </input>
<input>
<ID>IN_2</ID>594 </input>
<input>
<ID>IN_3</ID>599 </input>
<input>
<ID>IN_4</ID>598 </input>
<input>
<ID>IN_5</ID>593 </input>
<input>
<ID>IN_6</ID>596 </input>
<input>
<ID>IN_7</ID>595 </input>
<output>
<ID>OUT_0</ID>634 </output>
<output>
<ID>OUT_1</ID>635 </output>
<output>
<ID>OUT_2</ID>636 </output>
<output>
<ID>OUT_3</ID>637 </output>
<output>
<ID>OUT_4</ID>638 </output>
<output>
<ID>OUT_5</ID>639 </output>
<output>
<ID>OUT_6</ID>640 </output>
<output>
<ID>OUT_7</ID>641 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>111</ID>
<type>DA_FROM</type>
<position>18,-10.5</position>
<input>
<ID>IN_0</ID>189 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I3</lparam></gate>
<gate>
<ID>691</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>103,-44</position>
<input>
<ID>ENABLE_0</ID>605 </input>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>602 </input>
<input>
<ID>IN_2</ID>601 </input>
<input>
<ID>IN_3</ID>604 </input>
<output>
<ID>OUT_0</ID>619 </output>
<output>
<ID>OUT_1</ID>620 </output>
<output>
<ID>OUT_2</ID>621 </output>
<output>
<ID>OUT_3</ID>633 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>693</ID>
<type>DA_FROM</type>
<position>99,-26</position>
<input>
<ID>IN_0</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-BUS</lparam></gate>
<gate>
<ID>115</ID>
<type>FF_GND</type>
<position>35,-26.5</position>
<output>
<ID>OUT_0</ID>193 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>694</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>69.5,-54</position>
<input>
<ID>ENABLE_0</ID>618 </input>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>602 </input>
<input>
<ID>IN_2</ID>601 </input>
<input>
<ID>IN_3</ID>604 </input>
<output>
<ID>OUT_0</ID>606 </output>
<output>
<ID>OUT_1</ID>607 </output>
<output>
<ID>OUT_2</ID>608 </output>
<output>
<ID>OUT_3</ID>609 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>695</ID>
<type>DE_TO</type>
<position>67,-61</position>
<input>
<ID>IN_0</ID>606 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 0</lparam></gate>
<gate>
<ID>696</ID>
<type>DE_TO</type>
<position>69,-61</position>
<input>
<ID>IN_0</ID>607 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 1</lparam></gate>
<gate>
<ID>697</ID>
<type>DE_TO</type>
<position>71,-61</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 2</lparam></gate>
<gate>
<ID>698</ID>
<type>DE_TO</type>
<position>73,-61</position>
<input>
<ID>IN_0</ID>609 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 3</lparam></gate>
<gate>
<ID>699</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>78.5,-54</position>
<input>
<ID>ENABLE_0</ID>618 </input>
<input>
<ID>IN_0</ID>600 </input>
<input>
<ID>IN_1</ID>597 </input>
<input>
<ID>IN_2</ID>594 </input>
<input>
<ID>IN_3</ID>599 </input>
<output>
<ID>OUT_0</ID>610 </output>
<output>
<ID>OUT_1</ID>611 </output>
<output>
<ID>OUT_2</ID>612 </output>
<output>
<ID>OUT_3</ID>613 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>700</ID>
<type>DE_TO</type>
<position>76,-61</position>
<input>
<ID>IN_0</ID>610 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 4</lparam></gate>
<gate>
<ID>701</ID>
<type>DE_TO</type>
<position>78,-61</position>
<input>
<ID>IN_0</ID>611 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 5</lparam></gate>
<gate>
<ID>702</ID>
<type>DE_TO</type>
<position>80,-61</position>
<input>
<ID>IN_0</ID>612 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 6</lparam></gate>
<gate>
<ID>703</ID>
<type>DE_TO</type>
<position>82,-61</position>
<input>
<ID>IN_0</ID>613 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 7</lparam></gate>
<gate>
<ID>704</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>88,-54</position>
<input>
<ID>ENABLE_0</ID>618 </input>
<input>
<ID>IN_0</ID>598 </input>
<input>
<ID>IN_1</ID>593 </input>
<input>
<ID>IN_2</ID>596 </input>
<input>
<ID>IN_3</ID>595 </input>
<output>
<ID>OUT_0</ID>614 </output>
<output>
<ID>OUT_1</ID>615 </output>
<output>
<ID>OUT_2</ID>616 </output>
<output>
<ID>OUT_3</ID>617 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>705</ID>
<type>DE_TO</type>
<position>85.5,-61</position>
<input>
<ID>IN_0</ID>614 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 8</lparam></gate>
<gate>
<ID>706</ID>
<type>DE_TO</type>
<position>87.5,-61</position>
<input>
<ID>IN_0</ID>615 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 9</lparam></gate>
<gate>
<ID>707</ID>
<type>DE_TO</type>
<position>89.5,-61</position>
<input>
<ID>IN_0</ID>616 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 10</lparam></gate>
<gate>
<ID>708</ID>
<type>DE_TO</type>
<position>91.5,-61</position>
<input>
<ID>IN_0</ID>617 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 11</lparam></gate>
<gate>
<ID>709</ID>
<type>DA_FROM</type>
<position>96,-54</position>
<input>
<ID>IN_0</ID>618 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PC-ADDR</lparam></gate>
<gate>
<ID>710</ID>
<type>DE_TO</type>
<position>156,-48.5</position>
<input>
<ID>IN_0</ID>645 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>711</ID>
<type>DE_TO</type>
<position>152,-49</position>
<input>
<ID>IN_0</ID>644 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>712</ID>
<type>DE_TO</type>
<position>148.5,-49.5</position>
<input>
<ID>IN_0</ID>643 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>713</ID>
<type>DE_TO</type>
<position>145.5,-49.5</position>
<input>
<ID>IN_0</ID>642 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>714</ID>
<type>DE_TO</type>
<position>142,-49.5</position>
<input>
<ID>IN_0</ID>641 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>715</ID>
<type>DE_TO</type>
<position>138.5,-49.5</position>
<input>
<ID>IN_0</ID>640 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>716</ID>
<type>DE_TO</type>
<position>135.5,-50</position>
<input>
<ID>IN_0</ID>639 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>717</ID>
<type>DE_TO</type>
<position>132,-50</position>
<input>
<ID>IN_0</ID>638 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>718</ID>
<type>DE_TO</type>
<position>107.5,-50.5</position>
<input>
<ID>IN_0</ID>619 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>719</ID>
<type>DE_TO</type>
<position>111,-50.5</position>
<input>
<ID>IN_0</ID>620 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>720</ID>
<type>DE_TO</type>
<position>114,-50.5</position>
<input>
<ID>IN_0</ID>621 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>721</ID>
<type>DE_TO</type>
<position>117,-50.5</position>
<input>
<ID>IN_0</ID>633 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>722</ID>
<type>DE_TO</type>
<position>120,-50.5</position>
<input>
<ID>IN_0</ID>634 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>723</ID>
<type>DE_TO</type>
<position>122.5,-50.5</position>
<input>
<ID>IN_0</ID>635 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>724</ID>
<type>DE_TO</type>
<position>125,-50</position>
<input>
<ID>IN_0</ID>636 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>725</ID>
<type>DE_TO</type>
<position>128.5,-50</position>
<input>
<ID>IN_0</ID>637 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>727</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>112.5,-29</position>
<input>
<ID>ENABLE_0</ID>605 </input>
<input>
<ID>IN_0</ID>646 </input>
<input>
<ID>IN_1</ID>646 </input>
<input>
<ID>IN_2</ID>646 </input>
<input>
<ID>IN_3</ID>646 </input>
<output>
<ID>OUT_0</ID>642 </output>
<output>
<ID>OUT_1</ID>643 </output>
<output>
<ID>OUT_2</ID>644 </output>
<output>
<ID>OUT_3</ID>645 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>729</ID>
<type>FF_GND</type>
<position>109.5,-32.5</position>
<output>
<ID>OUT_0</ID>646 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>734</ID>
<type>DA_FROM</type>
<position>-77,3</position>
<input>
<ID>IN_0</ID>53 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>735</ID>
<type>DA_FROM</type>
<position>-77,5.5</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>736</ID>
<type>DA_FROM</type>
<position>-77,8</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>737</ID>
<type>DA_FROM</type>
<position>-77,10.5</position>
<input>
<ID>IN_0</ID>701 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>739</ID>
<type>AE_FULLADDER_4BIT</type>
<position>26,-27.5</position>
<input>
<ID>IN_0</ID>192 </input>
<input>
<ID>IN_1</ID>191 </input>
<input>
<ID>IN_2</ID>190 </input>
<input>
<ID>IN_3</ID>189 </input>
<input>
<ID>IN_B_0</ID>663 </input>
<input>
<ID>IN_B_1</ID>664 </input>
<input>
<ID>IN_B_2</ID>665 </input>
<input>
<ID>IN_B_3</ID>666 </input>
<output>
<ID>OUT_0</ID>649 </output>
<output>
<ID>OUT_1</ID>650 </output>
<output>
<ID>OUT_2</ID>651 </output>
<output>
<ID>OUT_3</ID>652 </output>
<input>
<ID>carry_in</ID>193 </input>
<output>
<ID>carry_out</ID>647 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>740</ID>
<type>AE_FULLADDER_4BIT</type>
<position>6,-27.5</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>187 </input>
<input>
<ID>IN_2</ID>186 </input>
<input>
<ID>IN_3</ID>184 </input>
<input>
<ID>IN_B_0</ID>671 </input>
<input>
<ID>IN_B_1</ID>672 </input>
<input>
<ID>IN_B_2</ID>673 </input>
<input>
<ID>IN_B_3</ID>674 </input>
<output>
<ID>OUT_0</ID>653 </output>
<output>
<ID>OUT_1</ID>654 </output>
<output>
<ID>OUT_2</ID>655 </output>
<output>
<ID>OUT_3</ID>656 </output>
<input>
<ID>carry_in</ID>647 </input>
<output>
<ID>carry_out</ID>648 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>741</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-15,-27.5</position>
<input>
<ID>IN_0</ID>180 </input>
<input>
<ID>IN_1</ID>181 </input>
<input>
<ID>IN_2</ID>182 </input>
<input>
<ID>IN_3</ID>183 </input>
<input>
<ID>IN_B_0</ID>676 </input>
<input>
<ID>IN_B_1</ID>677 </input>
<input>
<ID>IN_B_2</ID>678 </input>
<input>
<ID>IN_B_3</ID>679 </input>
<output>
<ID>OUT_0</ID>657 </output>
<output>
<ID>OUT_1</ID>658 </output>
<output>
<ID>OUT_2</ID>659 </output>
<output>
<ID>OUT_3</ID>660 </output>
<input>
<ID>carry_in</ID>648 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>747</ID>
<type>AA_AND2</type>
<position>51,-20</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>667 </input>
<output>
<ID>OUT</ID>663 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>748</ID>
<type>AA_AND2</type>
<position>50.5,-15</position>
<input>
<ID>IN_0</ID>602 </input>
<input>
<ID>IN_1</ID>667 </input>
<output>
<ID>OUT</ID>664 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>749</ID>
<type>AA_AND2</type>
<position>50.5,-10</position>
<input>
<ID>IN_0</ID>601 </input>
<input>
<ID>IN_1</ID>667 </input>
<output>
<ID>OUT</ID>665 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>750</ID>
<type>AA_AND2</type>
<position>50,-5</position>
<input>
<ID>IN_0</ID>604 </input>
<input>
<ID>IN_1</ID>667 </input>
<output>
<ID>OUT</ID>666 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>752</ID>
<type>DA_FROM</type>
<position>64.5,-4</position>
<input>
<ID>IN_0</ID>667 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Offset</lparam></gate>
<gate>
<ID>760</ID>
<type>AA_AND2</type>
<position>70,1.5</position>
<input>
<ID>IN_0</ID>600 </input>
<input>
<ID>IN_1</ID>670 </input>
<output>
<ID>OUT</ID>671 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>761</ID>
<type>AA_AND2</type>
<position>69.5,6.5</position>
<input>
<ID>IN_0</ID>597 </input>
<input>
<ID>IN_1</ID>670 </input>
<output>
<ID>OUT</ID>672 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>762</ID>
<type>AA_AND2</type>
<position>69.5,11.5</position>
<input>
<ID>IN_0</ID>594 </input>
<input>
<ID>IN_1</ID>670 </input>
<output>
<ID>OUT</ID>673 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>763</ID>
<type>AA_AND2</type>
<position>69,16.5</position>
<input>
<ID>IN_0</ID>599 </input>
<input>
<ID>IN_1</ID>670 </input>
<output>
<ID>OUT</ID>674 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>764</ID>
<type>DA_FROM</type>
<position>79.5,17.5</position>
<input>
<ID>IN_0</ID>670 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Offset</lparam></gate>
<gate>
<ID>765</ID>
<type>AA_AND2</type>
<position>79.5,24</position>
<input>
<ID>IN_0</ID>598 </input>
<input>
<ID>IN_1</ID>675 </input>
<output>
<ID>OUT</ID>676 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>766</ID>
<type>AA_AND2</type>
<position>79,29</position>
<input>
<ID>IN_0</ID>593 </input>
<input>
<ID>IN_1</ID>675 </input>
<output>
<ID>OUT</ID>677 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>767</ID>
<type>AA_AND2</type>
<position>79,34</position>
<input>
<ID>IN_0</ID>596 </input>
<input>
<ID>IN_1</ID>675 </input>
<output>
<ID>OUT</ID>678 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>768</ID>
<type>AA_AND2</type>
<position>78.5,39</position>
<input>
<ID>IN_0</ID>595 </input>
<input>
<ID>IN_1</ID>675 </input>
<output>
<ID>OUT</ID>679 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>769</ID>
<type>DA_FROM</type>
<position>93,40</position>
<input>
<ID>IN_0</ID>675 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Offset</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-26.5,34,-26.5</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<connection>
<GID>739</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-73,7.5,-73,8</points>
<intersection>7.5 1</intersection>
<intersection>8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-73,7.5,-71,7.5</points>
<connection>
<GID>812</GID>
<name>IN_2</name></connection>
<intersection>-73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75,8,-73,8</points>
<connection>
<GID>736</GID>
<name>IN_0</name></connection>
<intersection>-73 0</intersection></hsegment></shape></wire>
<wire>
<ID>588</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-49,53.5,-47</points>
<connection>
<GID>677</GID>
<name>clock</name></connection>
<connection>
<GID>679</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-51.5,55.5,-47</points>
<connection>
<GID>677</GID>
<name>clear</name></connection>
<connection>
<GID>681</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-32,55.5,-29.5</points>
<connection>
<GID>677</GID>
<name>count_up</name></connection>
<connection>
<GID>683</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-32,53.5,-30</points>
<connection>
<GID>677</GID>
<name>load</name></connection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-30,53.5,-30</points>
<connection>
<GID>685</GID>
<name>IN_0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-32,54.5,-24.5</points>
<connection>
<GID>677</GID>
<name>count_enable</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-24.5,54.5,-24.5</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-36,101,-36</points>
<connection>
<GID>677</GID>
<name>OUT_9</name></connection>
<connection>
<GID>689</GID>
<name>IN_5</name></connection>
<intersection>87.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>87.5,-52,87.5,28</points>
<connection>
<GID>704</GID>
<name>IN_1</name></connection>
<intersection>-36 1</intersection>
<intersection>28 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>82,28,87.5,28</points>
<connection>
<GID>766</GID>
<name>IN_0</name></connection>
<intersection>87.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-39,101,-39</points>
<connection>
<GID>677</GID>
<name>OUT_6</name></connection>
<connection>
<GID>689</GID>
<name>IN_2</name></connection>
<intersection>79 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>79,-52,79,10.5</points>
<connection>
<GID>699</GID>
<name>IN_2</name></connection>
<intersection>-39 1</intersection>
<intersection>10.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>72.5,10.5,79,10.5</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<intersection>79 3</intersection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-34,101,-34</points>
<connection>
<GID>677</GID>
<name>OUT_11</name></connection>
<connection>
<GID>689</GID>
<name>IN_7</name></connection>
<intersection>89.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>89.5,-52,89.5,38</points>
<connection>
<GID>704</GID>
<name>IN_3</name></connection>
<intersection>-34 1</intersection>
<intersection>38 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>81.5,38,89.5,38</points>
<connection>
<GID>768</GID>
<name>IN_0</name></connection>
<intersection>89.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-35,101,-35</points>
<connection>
<GID>677</GID>
<name>OUT_10</name></connection>
<connection>
<GID>689</GID>
<name>IN_6</name></connection>
<intersection>88.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>88.5,-52,88.5,33</points>
<connection>
<GID>704</GID>
<name>IN_2</name></connection>
<intersection>-35 1</intersection>
<intersection>33 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>82,33,88.5,33</points>
<connection>
<GID>767</GID>
<name>IN_0</name></connection>
<intersection>88.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-40,101,-40</points>
<connection>
<GID>677</GID>
<name>OUT_5</name></connection>
<connection>
<GID>689</GID>
<name>IN_1</name></connection>
<intersection>78 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>78,-52,78,5.5</points>
<connection>
<GID>699</GID>
<name>IN_1</name></connection>
<intersection>-40 1</intersection>
<intersection>5.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>72.5,5.5,78,5.5</points>
<connection>
<GID>761</GID>
<name>IN_0</name></connection>
<intersection>78 3</intersection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-37,101,-37</points>
<connection>
<GID>677</GID>
<name>OUT_8</name></connection>
<connection>
<GID>689</GID>
<name>IN_4</name></connection>
<intersection>86.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>86.5,-52,86.5,23</points>
<connection>
<GID>704</GID>
<name>IN_0</name></connection>
<intersection>-37 1</intersection>
<intersection>23 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>82.5,23,86.5,23</points>
<connection>
<GID>765</GID>
<name>IN_0</name></connection>
<intersection>86.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-38,101,-38</points>
<connection>
<GID>677</GID>
<name>OUT_7</name></connection>
<connection>
<GID>689</GID>
<name>IN_3</name></connection>
<intersection>80 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>80,-52,80,15.5</points>
<connection>
<GID>699</GID>
<name>IN_3</name></connection>
<intersection>-38 1</intersection>
<intersection>15.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>72,15.5,80,15.5</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<intersection>80 3</intersection></hsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-41,101,-41</points>
<connection>
<GID>677</GID>
<name>OUT_4</name></connection>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<intersection>77 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77,-52,77,0.5</points>
<connection>
<GID>699</GID>
<name>IN_0</name></connection>
<intersection>-41 1</intersection>
<intersection>0.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>73,0.5,77,0.5</points>
<connection>
<GID>760</GID>
<name>IN_0</name></connection>
<intersection>77 3</intersection></hsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-43.5,101,-43.5</points>
<connection>
<GID>691</GID>
<name>IN_2</name></connection>
<intersection>70 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>70,-52,70,-11</points>
<connection>
<GID>694</GID>
<name>IN_2</name></connection>
<intersection>-43.5 1</intersection>
<intersection>-43 9</intersection>
<intersection>-11 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>53.5,-11,70,-11</points>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<intersection>70 5</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>59.5,-43,70,-43</points>
<connection>
<GID>677</GID>
<name>OUT_2</name></connection>
<intersection>70 5</intersection></hsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,-44.5,101,-44.5</points>
<connection>
<GID>691</GID>
<name>IN_1</name></connection>
<intersection>69 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>69,-52,69,-16</points>
<connection>
<GID>694</GID>
<name>IN_1</name></connection>
<intersection>-44.5 1</intersection>
<intersection>-44 13</intersection>
<intersection>-16 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>53.5,-16,69,-16</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<intersection>69 5</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>59.5,-44,69,-44</points>
<connection>
<GID>677</GID>
<name>OUT_1</name></connection>
<intersection>69 5</intersection></hsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-45.5,101,-45.5</points>
<connection>
<GID>691</GID>
<name>IN_0</name></connection>
<intersection>68 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>68,-52,68,-21</points>
<connection>
<GID>694</GID>
<name>IN_0</name></connection>
<intersection>-45.5 1</intersection>
<intersection>-45 11</intersection>
<intersection>-21 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>54,-21,68,-21</points>
<connection>
<GID>747</GID>
<name>IN_0</name></connection>
<intersection>68 5</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>59.5,-45,68,-45</points>
<connection>
<GID>677</GID>
<name>OUT_0</name></connection>
<intersection>68 5</intersection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-42,100.5,-42</points>
<connection>
<GID>677</GID>
<name>OUT_3</name></connection>
<intersection>71 5</intersection>
<intersection>100.5 7</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>71,-52,71,-6</points>
<connection>
<GID>694</GID>
<name>IN_3</name></connection>
<intersection>-42 1</intersection>
<intersection>-6 10</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>100.5,-42.5,100.5,-42</points>
<intersection>-42.5 8</intersection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>100.5,-42.5,101,-42.5</points>
<connection>
<GID>691</GID>
<name>IN_3</name></connection>
<intersection>100.5 7</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>53,-6,71,-6</points>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<intersection>71 5</intersection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-41,103,-26</points>
<connection>
<GID>689</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>691</GID>
<name>ENABLE_0</name></connection>
<intersection>-26 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>101,-26,112.5,-26</points>
<connection>
<GID>727</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>693</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-59,67,-56</points>
<connection>
<GID>695</GID>
<name>IN_0</name></connection>
<intersection>-56 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>67,-56,68,-56</points>
<connection>
<GID>694</GID>
<name>OUT_0</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-59,69,-56</points>
<connection>
<GID>696</GID>
<name>IN_0</name></connection>
<connection>
<GID>694</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-59,71,-56</points>
<connection>
<GID>697</GID>
<name>IN_0</name></connection>
<intersection>-56 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-56,71,-56</points>
<connection>
<GID>694</GID>
<name>OUT_2</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-56.5,71,-56</points>
<connection>
<GID>694</GID>
<name>OUT_3</name></connection>
<intersection>-56.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>73,-59,73,-56.5</points>
<connection>
<GID>698</GID>
<name>IN_0</name></connection>
<intersection>-56.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>71,-56.5,73,-56.5</points>
<intersection>71 0</intersection>
<intersection>73 1</intersection></hsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-59,76,-56</points>
<connection>
<GID>700</GID>
<name>IN_0</name></connection>
<intersection>-56 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>76,-56,77,-56</points>
<connection>
<GID>699</GID>
<name>OUT_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-59,78,-56</points>
<connection>
<GID>701</GID>
<name>IN_0</name></connection>
<connection>
<GID>699</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-59,80,-57.5</points>
<connection>
<GID>702</GID>
<name>IN_0</name></connection>
<intersection>-57.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-57.5,80,-57.5</points>
<intersection>79 5</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>79,-57.5,79,-56</points>
<connection>
<GID>699</GID>
<name>OUT_2</name></connection>
<intersection>-57.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>82,-59,82,-56</points>
<connection>
<GID>703</GID>
<name>IN_0</name></connection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>80,-56,82,-56</points>
<connection>
<GID>699</GID>
<name>OUT_3</name></connection>
<intersection>82 1</intersection></hsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-59,85.5,-56</points>
<connection>
<GID>705</GID>
<name>IN_0</name></connection>
<intersection>-56 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>85.5,-56,86.5,-56</points>
<connection>
<GID>704</GID>
<name>OUT_0</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-59,87.5,-56</points>
<connection>
<GID>706</GID>
<name>IN_0</name></connection>
<connection>
<GID>704</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-59,89.5,-56</points>
<connection>
<GID>707</GID>
<name>IN_0</name></connection>
<intersection>-56 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>88.5,-56,89.5,-56</points>
<connection>
<GID>704</GID>
<name>OUT_2</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-56.5,89.5,-56</points>
<connection>
<GID>704</GID>
<name>OUT_3</name></connection>
<intersection>-56.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>91.5,-59,91.5,-56.5</points>
<connection>
<GID>708</GID>
<name>IN_0</name></connection>
<intersection>-56.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-56.5,91.5,-56.5</points>
<intersection>89.5 0</intersection>
<intersection>91.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72.5,-54,94,-54</points>
<connection>
<GID>704</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>699</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>694</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>709</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-48.5,107.5,-45.5</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-45.5,107.5,-45.5</points>
<connection>
<GID>691</GID>
<name>OUT_0</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-48.5,111,-44.5</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-44.5,111,-44.5</points>
<connection>
<GID>691</GID>
<name>OUT_1</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-48.5,114,-43.5</points>
<connection>
<GID>720</GID>
<name>IN_0</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-43.5,114,-43.5</points>
<connection>
<GID>691</GID>
<name>OUT_2</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-73,5.5,-73,6.5</points>
<intersection>5.5 2</intersection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-73,6.5,-71,6.5</points>
<connection>
<GID>812</GID>
<name>IN_1</name></connection>
<intersection>-73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75,5.5,-73,5.5</points>
<connection>
<GID>735</GID>
<name>IN_0</name></connection>
<intersection>-73 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72,3,-72,5.5</points>
<intersection>3 2</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72,5.5,-71,5.5</points>
<connection>
<GID>812</GID>
<name>IN_0</name></connection>
<intersection>-72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75,3,-72,3</points>
<connection>
<GID>734</GID>
<name>IN_0</name></connection>
<intersection>-72 0</intersection></hsegment></shape></wire>
<wire>
<ID>633</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,-48.5,117,-42.5</points>
<connection>
<GID>721</GID>
<name>IN_0</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-42.5,117,-42.5</points>
<connection>
<GID>691</GID>
<name>OUT_3</name></connection>
<intersection>117 0</intersection></hsegment></shape></wire>
<wire>
<ID>634</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-48.5,120,-41</points>
<connection>
<GID>722</GID>
<name>IN_0</name></connection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-41,120,-41</points>
<connection>
<GID>689</GID>
<name>OUT_0</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>635</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-48.5,122.5,-40</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-40,122.5,-40</points>
<connection>
<GID>689</GID>
<name>OUT_1</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7,-57.5,-3,-57.5</points>
<connection>
<GID>275</GID>
<name>OUT_0</name></connection>
<connection>
<GID>276</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>636</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-48,125,-39</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-39,125,-39</points>
<connection>
<GID>689</GID>
<name>OUT_2</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-48,128.5,-38</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-38,128.5,-38</points>
<connection>
<GID>689</GID>
<name>OUT_3</name></connection>
<intersection>128.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>638</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-48,132,-37</points>
<connection>
<GID>717</GID>
<name>IN_0</name></connection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-37,132,-37</points>
<connection>
<GID>689</GID>
<name>OUT_4</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>639</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-48,135.5,-36</points>
<connection>
<GID>716</GID>
<name>IN_0</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-36,135.5,-36</points>
<connection>
<GID>689</GID>
<name>OUT_5</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-47.5,138.5,-35</points>
<connection>
<GID>715</GID>
<name>IN_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-35,138.5,-35</points>
<connection>
<GID>689</GID>
<name>OUT_6</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>641</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-47.5,142,-34</points>
<connection>
<GID>714</GID>
<name>IN_0</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-34,142,-34</points>
<connection>
<GID>689</GID>
<name>OUT_7</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>642</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-47.5,145.5,-30.5</points>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-30.5,145.5,-30.5</points>
<connection>
<GID>727</GID>
<name>OUT_0</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-47.5,148.5,-29.5</points>
<connection>
<GID>712</GID>
<name>IN_0</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-29.5,148.5,-29.5</points>
<connection>
<GID>727</GID>
<name>OUT_1</name></connection>
<intersection>148.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>644</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,-47,152,-28.5</points>
<connection>
<GID>711</GID>
<name>IN_0</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-28.5,152,-28.5</points>
<connection>
<GID>727</GID>
<name>OUT_2</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>645</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-46.5,156,-27.5</points>
<connection>
<GID>710</GID>
<name>IN_0</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-27.5,156,-27.5</points>
<connection>
<GID>727</GID>
<name>OUT_3</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>646</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-31.5,109.5,-30.5</points>
<connection>
<GID>729</GID>
<name>OUT_0</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-30.5,110.5,-30.5</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-30.5,110.5,-27.5</points>
<connection>
<GID>727</GID>
<name>IN_3</name></connection>
<connection>
<GID>727</GID>
<name>IN_2</name></connection>
<connection>
<GID>727</GID>
<name>IN_1</name></connection>
<intersection>-30.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-26.5,18,-26.5</points>
<connection>
<GID>739</GID>
<name>carry_out</name></connection>
<connection>
<GID>740</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7,-26.5,-2,-26.5</points>
<connection>
<GID>740</GID>
<name>carry_out</name></connection>
<connection>
<GID>741</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-45,27.5,-31.5</points>
<connection>
<GID>739</GID>
<name>OUT_0</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-45,49.5,-45</points>
<connection>
<GID>677</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-44,26.5,-31.5</points>
<connection>
<GID>739</GID>
<name>OUT_1</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-44,49.5,-44</points>
<connection>
<GID>677</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-43,25.5,-31.5</points>
<connection>
<GID>739</GID>
<name>OUT_2</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-43,49.5,-43</points>
<connection>
<GID>677</GID>
<name>IN_2</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-42,24.5,-31.5</points>
<connection>
<GID>739</GID>
<name>OUT_3</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-42,49.5,-42</points>
<connection>
<GID>677</GID>
<name>IN_3</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>653</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-41,7.5,-31.5</points>
<connection>
<GID>740</GID>
<name>OUT_0</name></connection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,-41,49.5,-41</points>
<connection>
<GID>677</GID>
<name>IN_4</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>654</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-40,6.5,-31.5</points>
<connection>
<GID>740</GID>
<name>OUT_1</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-40,49.5,-40</points>
<connection>
<GID>677</GID>
<name>IN_5</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>655</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-39,5.5,-31.5</points>
<connection>
<GID>740</GID>
<name>OUT_2</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,-39,49.5,-39</points>
<connection>
<GID>677</GID>
<name>IN_6</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>656</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-38,4.5,-31.5</points>
<connection>
<GID>740</GID>
<name>OUT_3</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4.5,-38,49.5,-38</points>
<connection>
<GID>677</GID>
<name>IN_7</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>657</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-37,-13.5,-31.5</points>
<connection>
<GID>741</GID>
<name>OUT_0</name></connection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13.5,-37,49.5,-37</points>
<connection>
<GID>677</GID>
<name>IN_8</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-73,-1.5,-73,-1</points>
<intersection>-1.5 2</intersection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-75,-1,-73,-1</points>
<connection>
<GID>803</GID>
<name>IN_0</name></connection>
<intersection>-73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-73,-1.5,-67,-1.5</points>
<connection>
<GID>3</GID>
<name>IN_7</name></connection>
<intersection>-73 0</intersection></hsegment></shape></wire>
<wire>
<ID>658</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-36,-14.5,-31.5</points>
<connection>
<GID>741</GID>
<name>OUT_1</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-36,49.5,-36</points>
<connection>
<GID>677</GID>
<name>IN_9</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-73.5,-3.5,-73.5,-2.5</points>
<intersection>-3.5 1</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-74.5,-3.5,-73.5,-3.5</points>
<connection>
<GID>804</GID>
<name>IN_0</name></connection>
<intersection>-73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-73.5,-2.5,-67,-2.5</points>
<connection>
<GID>3</GID>
<name>IN_6</name></connection>
<intersection>-73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>659</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-35,-15.5,-31.5</points>
<connection>
<GID>741</GID>
<name>OUT_2</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15.5,-35,49.5,-35</points>
<connection>
<GID>677</GID>
<name>IN_10</name></connection>
<intersection>-15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-73,-6.5,-73,-3.5</points>
<intersection>-6.5 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-75.5,-6.5,-73,-6.5</points>
<connection>
<GID>805</GID>
<name>IN_0</name></connection>
<intersection>-73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-73,-3.5,-67,-3.5</points>
<connection>
<GID>3</GID>
<name>IN_5</name></connection>
<intersection>-73 0</intersection></hsegment></shape></wire>
<wire>
<ID>660</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-34,-16.5,-31.5</points>
<connection>
<GID>741</GID>
<name>OUT_3</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16.5,-34,49.5,-34</points>
<connection>
<GID>677</GID>
<name>IN_11</name></connection>
<intersection>-16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71.5,-9.5,-71.5,-4.5</points>
<intersection>-9.5 1</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-74.5,-9.5,-71.5,-9.5</points>
<connection>
<GID>806</GID>
<name>IN_0</name></connection>
<intersection>-71.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-4.5,-67,-4.5</points>
<connection>
<GID>3</GID>
<name>IN_4</name></connection>
<intersection>-71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71,-11.5,-71,-5.5</points>
<intersection>-11.5 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-74.5,-11.5,-71,-11.5</points>
<connection>
<GID>807</GID>
<name>IN_0</name></connection>
<intersection>-71 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71,-5.5,-67,-5.5</points>
<connection>
<GID>3</GID>
<name>IN_3</name></connection>
<intersection>-71 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70.5,-14.5,-70.5,-6.5</points>
<intersection>-14.5 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-70.5,-6.5,-67,-6.5</points>
<connection>
<GID>3</GID>
<name>IN_2</name></connection>
<intersection>-70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-74.5,-14.5,-70.5,-14.5</points>
<connection>
<GID>808</GID>
<name>IN_0</name></connection>
<intersection>-70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-23.5,31,-20</points>
<connection>
<GID>739</GID>
<name>IN_B_0</name></connection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-20,48,-20</points>
<connection>
<GID>747</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69.5,-17.5,-69.5,-7.5</points>
<intersection>-17.5 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,-7.5,-67,-7.5</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>-69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75,-17.5,-69.5,-17.5</points>
<connection>
<GID>809</GID>
<name>IN_0</name></connection>
<intersection>-69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>664</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-23.5,30,-15</points>
<connection>
<GID>739</GID>
<name>IN_B_1</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-15,47.5,-15</points>
<connection>
<GID>748</GID>
<name>OUT</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68.5,-21.5,-68.5,-8.5</points>
<intersection>-21.5 1</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-75,-21.5,-68.5,-21.5</points>
<connection>
<GID>810</GID>
<name>IN_0</name></connection>
<intersection>-68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-68.5,-8.5,-67,-8.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>-68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>665</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-23.5,29,-10</points>
<connection>
<GID>739</GID>
<name>IN_B_2</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-10,47.5,-10</points>
<connection>
<GID>749</GID>
<name>OUT</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-67,8.5,-62.5,8.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<connection>
<GID>812</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-23.5,28,-5</points>
<connection>
<GID>739</GID>
<name>IN_B_3</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-5,47,-5</points>
<connection>
<GID>750</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64,6.5,-64,7.5</points>
<intersection>6.5 2</intersection>
<intersection>7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67,7.5,-64,7.5</points>
<connection>
<GID>812</GID>
<name>OUT_2</name></connection>
<intersection>-64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-64,6.5,-62.5,6.5</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>-64 0</intersection></hsegment></shape></wire>
<wire>
<ID>667</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>53,-4,62.5,-4</points>
<connection>
<GID>750</GID>
<name>IN_1</name></connection>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<intersection>54.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54.5,-19,54.5,-4</points>
<intersection>-19 8</intersection>
<intersection>-14 5</intersection>
<intersection>-9 6</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>53.5,-14,54.5,-14</points>
<connection>
<GID>748</GID>
<name>IN_1</name></connection>
<intersection>54.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>53.5,-9,54.5,-9</points>
<connection>
<GID>749</GID>
<name>IN_1</name></connection>
<intersection>54.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>54,-19,54.5,-19</points>
<connection>
<GID>747</GID>
<name>IN_1</name></connection>
<intersection>54.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,4,-64.5,6.5</points>
<intersection>4 2</intersection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67,6.5,-64.5,6.5</points>
<connection>
<GID>812</GID>
<name>OUT_1</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-64.5,4,-62.5,4</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,2,-65,5.5</points>
<intersection>2 2</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67,5.5,-65,5.5</points>
<connection>
<GID>812</GID>
<name>OUT_0</name></connection>
<intersection>-65 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-65,2,-62.5,2</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-65 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-63,-1.5,-51.5,-1.5</points>
<connection>
<GID>3</GID>
<name>OUT_7</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>670</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>72,17.5,77.5,17.5</points>
<connection>
<GID>763</GID>
<name>IN_1</name></connection>
<connection>
<GID>764</GID>
<name>IN_0</name></connection>
<intersection>73.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>73.5,2.5,73.5,17.5</points>
<intersection>2.5 8</intersection>
<intersection>7.5 5</intersection>
<intersection>12.5 6</intersection>
<intersection>17.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>72.5,7.5,73.5,7.5</points>
<connection>
<GID>761</GID>
<name>IN_1</name></connection>
<intersection>73.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>72.5,12.5,73.5,12.5</points>
<connection>
<GID>762</GID>
<name>IN_1</name></connection>
<intersection>73.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>73,2.5,73.5,2.5</points>
<connection>
<GID>760</GID>
<name>IN_1</name></connection>
<intersection>73.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52.5,-3.5,-52.5,-2.5</points>
<intersection>-3.5 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63,-2.5,-52.5,-2.5</points>
<connection>
<GID>3</GID>
<name>OUT_6</name></connection>
<intersection>-52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,-3.5,-51.5,-3.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>-52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>671</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-23.5,11,1.5</points>
<connection>
<GID>740</GID>
<name>IN_B_0</name></connection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,1.5,67,1.5</points>
<connection>
<GID>760</GID>
<name>OUT</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53.5,-6,-53.5,-3.5</points>
<intersection>-6 2</intersection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63,-3.5,-53.5,-3.5</points>
<connection>
<GID>3</GID>
<name>OUT_5</name></connection>
<intersection>-53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-53.5,-6,-51.5,-6</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-23.5,10,6.5</points>
<connection>
<GID>740</GID>
<name>IN_B_1</name></connection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,6.5,66.5,6.5</points>
<connection>
<GID>761</GID>
<name>OUT</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54.5,-8,-54.5,-4.5</points>
<intersection>-8 1</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54.5,-8,-51.5,-8</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-63,-4.5,-54.5,-4.5</points>
<connection>
<GID>3</GID>
<name>OUT_4</name></connection>
<intersection>-54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>673</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-23.5,9,11.5</points>
<connection>
<GID>740</GID>
<name>IN_B_2</name></connection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,11.5,66.5,11.5</points>
<connection>
<GID>762</GID>
<name>OUT</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-23.5,8,16.5</points>
<connection>
<GID>740</GID>
<name>IN_B_3</name></connection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,16.5,66,16.5</points>
<connection>
<GID>763</GID>
<name>OUT</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>675</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>81.5,40,91,40</points>
<connection>
<GID>768</GID>
<name>IN_1</name></connection>
<connection>
<GID>769</GID>
<name>IN_0</name></connection>
<intersection>83 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>83,25,83,40</points>
<intersection>25 8</intersection>
<intersection>30 5</intersection>
<intersection>35 6</intersection>
<intersection>40 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>82,30,83,30</points>
<connection>
<GID>766</GID>
<name>IN_1</name></connection>
<intersection>83 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>82,35,83,35</points>
<connection>
<GID>767</GID>
<name>IN_1</name></connection>
<intersection>83 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>82.5,25,83,25</points>
<connection>
<GID>765</GID>
<name>IN_1</name></connection>
<intersection>83 3</intersection></hsegment></shape></wire>
<wire>
<ID>676</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-23.5,-10,24</points>
<connection>
<GID>741</GID>
<name>IN_B_0</name></connection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,24,76.5,24</points>
<connection>
<GID>765</GID>
<name>OUT</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>677</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-23.5,-11,29</points>
<connection>
<GID>741</GID>
<name>IN_B_1</name></connection>
<intersection>29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11,29,76,29</points>
<connection>
<GID>766</GID>
<name>OUT</name></connection>
<intersection>-11 0</intersection></hsegment></shape></wire>
<wire>
<ID>678</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-23.5,-12,34</points>
<connection>
<GID>741</GID>
<name>IN_B_2</name></connection>
<intersection>34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,34,76,34</points>
<connection>
<GID>767</GID>
<name>OUT</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-23.5,-13,39</points>
<connection>
<GID>741</GID>
<name>IN_B_3</name></connection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,39,75.5,39</points>
<connection>
<GID>768</GID>
<name>OUT</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-73,8.5,-73,10.5</points>
<intersection>8.5 2</intersection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-75,10.5,-73,10.5</points>
<connection>
<GID>737</GID>
<name>IN_0</name></connection>
<intersection>-73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-73,8.5,-71,8.5</points>
<connection>
<GID>812</GID>
<name>IN_3</name></connection>
<intersection>-73 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,-10.5,-57.5,-5.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-63,-5.5,-57.5,-5.5</points>
<connection>
<GID>3</GID>
<name>OUT_3</name></connection>
<intersection>-57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58.5,-12.5,-58.5,-6.5</points>
<intersection>-12.5 1</intersection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58.5,-12.5,-57.5,-12.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-63,-6.5,-58.5,-6.5</points>
<connection>
<GID>3</GID>
<name>OUT_2</name></connection>
<intersection>-58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59.5,-15,-59.5,-7.5</points>
<intersection>-15 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59.5,-15,-57.5,-15</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-63,-7.5,-59.5,-7.5</points>
<connection>
<GID>3</GID>
<name>OUT_1</name></connection>
<intersection>-59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60.5,-17,-60.5,-8.5</points>
<intersection>-17 1</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60.5,-17,-57.5,-17</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>-60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-63,-8.5,-60.5,-8.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69,0,-69,20.5</points>
<connection>
<GID>812</GID>
<name>ENABLE_0</name></connection>
<intersection>0 2</intersection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-79.5,20.5,-69,20.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69,0,-65,0</points>
<connection>
<GID>3</GID>
<name>ENABLE_0</name></connection>
<intersection>-69 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,-23.5,-17,-18</points>
<connection>
<GID>741</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-15.5,-18,-15.5,-12.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-17,-18,-15.5,-18</points>
<intersection>-17 0</intersection>
<intersection>-15.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18,-23.5,-18,-12.5</points>
<connection>
<GID>741</GID>
<name>IN_1</name></connection>
<connection>
<GID>61</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19,-23.5,-19,-18</points>
<connection>
<GID>741</GID>
<name>IN_2</name></connection>
<intersection>-18 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-20.5,-18,-20.5,-12.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-20.5,-18,-19,-18</points>
<intersection>-20.5 1</intersection>
<intersection>-19 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,-23.5,-20,-19</points>
<connection>
<GID>741</GID>
<name>IN_3</name></connection>
<intersection>-19 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-23,-19,-23,-12.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-23,-19,-20,-19</points>
<intersection>-23 1</intersection>
<intersection>-20 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-23.5,1,-22</points>
<connection>
<GID>740</GID>
<name>IN_3</name></connection>
<intersection>-22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-2.5,-22,-2.5,-13</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-2.5,-22,1,-22</points>
<intersection>-2.5 1</intersection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-23.5,2,-21</points>
<connection>
<GID>740</GID>
<name>IN_2</name></connection>
<intersection>-21 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-7.30078e-008,-21,-7.30078e-008,-13</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-7.30078e-008,-21,2,-21</points>
<intersection>-7.30078e-008 1</intersection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-23.5,3,-18</points>
<connection>
<GID>740</GID>
<name>IN_1</name></connection>
<intersection>-18 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>2.5,-18,2.5,-13</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>2.5,-18,3,-18</points>
<intersection>2.5 1</intersection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-23.5,4,-18</points>
<connection>
<GID>740</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>5,-18,5,-13</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>4,-18,5,-18</points>
<intersection>4 0</intersection>
<intersection>5 1</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-23.5,21,-20.5</points>
<connection>
<GID>739</GID>
<name>IN_3</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>18,-20.5,18,-12.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>18,-20.5,21,-20.5</points>
<intersection>18 1</intersection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-23.5,22,-18</points>
<connection>
<GID>739</GID>
<name>IN_2</name></connection>
<intersection>-18 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>20.5,-18,20.5,-12.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-18,22,-18</points>
<intersection>20.5 1</intersection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-23.5,23,-12.5</points>
<connection>
<GID>739</GID>
<name>IN_1</name></connection>
<connection>
<GID>91</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-23.5,24,-18</points>
<connection>
<GID>739</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>25.5,-18,25.5,-12.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>24,-18,25.5,-18</points>
<intersection>24 0</intersection>
<intersection>25.5 1</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>400.186,136.146,1073.59,-250.195</PageViewport>
<gate>
<ID>203</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>509,66</position>
<input>
<ID>ENABLE_0</ID>628 </input>
<input>
<ID>IN_0</ID>622 </input>
<input>
<ID>IN_1</ID>582 </input>
<input>
<ID>IN_2</ID>581 </input>
<input>
<ID>IN_3</ID>623 </input>
<output>
<ID>OUT_0</ID>744 </output>
<output>
<ID>OUT_1</ID>745 </output>
<output>
<ID>OUT_2</ID>746 </output>
<output>
<ID>OUT_3</ID>747 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>791</ID>
<type>DA_FROM</type>
<position>439,61.5</position>
<input>
<ID>IN_0</ID>796 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>795</ID>
<type>DA_FROM</type>
<position>438.5,58.5</position>
<input>
<ID>IN_0</ID>786 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>796</ID>
<type>DA_FROM</type>
<position>438.5,55.5</position>
<input>
<ID>IN_0</ID>785 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>798</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>456.5,68</position>
<input>
<ID>ENABLE_0</ID>802 </input>
<input>
<ID>IN_0</ID>785 </input>
<input>
<ID>IN_1</ID>786 </input>
<input>
<ID>IN_2</ID>796 </input>
<input>
<ID>IN_3</ID>797 </input>
<input>
<ID>IN_4</ID>798 </input>
<input>
<ID>IN_5</ID>799 </input>
<input>
<ID>IN_6</ID>800 </input>
<input>
<ID>IN_7</ID>801 </input>
<output>
<ID>OUT_0</ID>780 </output>
<output>
<ID>OUT_1</ID>775 </output>
<output>
<ID>OUT_2</ID>776 </output>
<output>
<ID>OUT_3</ID>777 </output>
<output>
<ID>OUT_4</ID>778 </output>
<output>
<ID>OUT_5</ID>779 </output>
<output>
<ID>OUT_6</ID>774 </output>
<output>
<ID>OUT_7</ID>773 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>412</ID>
<type>DA_FROM</type>
<position>512,50.5</position>
<input>
<ID>IN_0</ID>729 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID ADREG-ADDR</lparam></gate>
<gate>
<ID>413</ID>
<type>DE_TO</type>
<position>554.5,61.5</position>
<input>
<ID>IN_0</ID>759 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>800</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>452.5,74</position>
<input>
<ID>ENABLE_0</ID>802 </input>
<input>
<ID>IN_0</ID>795 </input>
<input>
<ID>IN_1</ID>794 </input>
<input>
<ID>IN_2</ID>793 </input>
<input>
<ID>IN_3</ID>792 </input>
<output>
<ID>OUT_0</ID>782 </output>
<output>
<ID>OUT_1</ID>781 </output>
<output>
<ID>OUT_2</ID>784 </output>
<output>
<ID>OUT_3</ID>783 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>607</ID>
<type>DE_TO</type>
<position>518.5,61.5</position>
<input>
<ID>IN_0</ID>746 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>802</ID>
<type>DA_FROM</type>
<position>457.5,80.5</position>
<input>
<ID>IN_0</ID>802 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID BUS-ADREG</lparam></gate>
<gate>
<ID>609</ID>
<type>DE_TO</type>
<position>521.5,61.5</position>
<input>
<ID>IN_0</ID>747 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>811</ID>
<type>DA_FROM</type>
<position>430.5,24.5</position>
<input>
<ID>IN_0</ID>809 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>813</ID>
<type>DA_FROM</type>
<position>430,21.5</position>
<input>
<ID>IN_0</ID>804 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>620</ID>
<type>DE_TO</type>
<position>524.5,61.5</position>
<input>
<ID>IN_0</ID>748 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>814</ID>
<type>DA_FROM</type>
<position>430,18.5</position>
<input>
<ID>IN_0</ID>803 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>815</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>449.5,31</position>
<input>
<ID>ENABLE_0</ID>815 </input>
<input>
<ID>IN_0</ID>803 </input>
<input>
<ID>IN_1</ID>804 </input>
<input>
<ID>IN_2</ID>809 </input>
<input>
<ID>IN_3</ID>810 </input>
<input>
<ID>IN_4</ID>811 </input>
<input>
<ID>IN_5</ID>812 </input>
<input>
<ID>IN_6</ID>813 </input>
<input>
<ID>IN_7</ID>814 </input>
<output>
<ID>OUT_0</ID>780 </output>
<output>
<ID>OUT_1</ID>775 </output>
<output>
<ID>OUT_2</ID>776 </output>
<output>
<ID>OUT_3</ID>777 </output>
<output>
<ID>OUT_4</ID>778 </output>
<output>
<ID>OUT_5</ID>779 </output>
<output>
<ID>OUT_6</ID>774 </output>
<output>
<ID>OUT_7</ID>773 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>816</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>445,37</position>
<input>
<ID>ENABLE_0</ID>815 </input>
<input>
<ID>IN_0</ID>808 </input>
<input>
<ID>IN_1</ID>807 </input>
<input>
<ID>IN_2</ID>806 </input>
<input>
<ID>IN_3</ID>805 </input>
<output>
<ID>OUT_0</ID>782 </output>
<output>
<ID>OUT_1</ID>781 </output>
<output>
<ID>OUT_2</ID>784 </output>
<output>
<ID>OUT_3</ID>783 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>817</ID>
<type>DA_FROM</type>
<position>474,40</position>
<input>
<ID>IN_0</ID>815 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID RES-ADREG</lparam></gate>
<gate>
<ID>818</ID>
<type>DA_FROM</type>
<position>430.5,49</position>
<input>
<ID>IN_0</ID>805 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A11</lparam></gate>
<gate>
<ID>819</ID>
<type>DA_FROM</type>
<position>430.5,46</position>
<input>
<ID>IN_0</ID>806 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A10</lparam></gate>
<gate>
<ID>820</ID>
<type>DA_FROM</type>
<position>430.5,43.5</position>
<input>
<ID>IN_0</ID>807 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A9</lparam></gate>
<gate>
<ID>821</ID>
<type>DA_FROM</type>
<position>430.5,41</position>
<input>
<ID>IN_0</ID>808 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A8</lparam></gate>
<gate>
<ID>823</ID>
<type>DA_FROM</type>
<position>430.5,38</position>
<input>
<ID>IN_0</ID>814 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A7</lparam></gate>
<gate>
<ID>824</ID>
<type>DA_FROM</type>
<position>430.5,35.5</position>
<input>
<ID>IN_0</ID>813 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A6</lparam></gate>
<gate>
<ID>825</ID>
<type>DA_FROM</type>
<position>430.5,32.5</position>
<input>
<ID>IN_0</ID>812 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A5</lparam></gate>
<gate>
<ID>632</ID>
<type>DE_TO</type>
<position>527,61.5</position>
<input>
<ID>IN_0</ID>749 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>826</ID>
<type>DA_FROM</type>
<position>430.5,30</position>
<input>
<ID>IN_0</ID>811 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A4</lparam></gate>
<gate>
<ID>827</ID>
<type>DA_FROM</type>
<position>430.5,27.5</position>
<input>
<ID>IN_0</ID>810 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>263</ID>
<type>DA_FROM</type>
<position>507,84</position>
<input>
<ID>IN_0</ID>628 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADREG-BUS</lparam></gate>
<gate>
<ID>265</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>482.5,58</position>
<input>
<ID>ENABLE_0</ID>729 </input>
<input>
<ID>IN_0</ID>622 </input>
<input>
<ID>IN_1</ID>582 </input>
<input>
<ID>IN_2</ID>581 </input>
<input>
<ID>IN_3</ID>623 </input>
<output>
<ID>OUT_0</ID>714 </output>
<output>
<ID>OUT_1</ID>715 </output>
<output>
<ID>OUT_2</ID>716 </output>
<output>
<ID>OUT_3</ID>717 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>653</ID>
<type>DE_TO</type>
<position>529.5,62</position>
<input>
<ID>IN_0</ID>750 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>267</ID>
<type>DE_TO</type>
<position>479.5,51</position>
<input>
<ID>IN_0</ID>714 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 0</lparam></gate>
<gate>
<ID>654</ID>
<type>DE_TO</type>
<position>531.5,62</position>
<input>
<ID>IN_0</ID>751 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>655</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>519.5,81</position>
<input>
<ID>ENABLE_0</ID>628 </input>
<input>
<ID>IN_0</ID>760 </input>
<input>
<ID>IN_1</ID>760 </input>
<input>
<ID>IN_2</ID>760 </input>
<input>
<ID>IN_3</ID>760 </input>
<output>
<ID>OUT_0</ID>756 </output>
<output>
<ID>OUT_1</ID>757 </output>
<output>
<ID>OUT_2</ID>758 </output>
<output>
<ID>OUT_3</ID>759 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>269</ID>
<type>DE_TO</type>
<position>482,51</position>
<input>
<ID>IN_0</ID>715 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 1</lparam></gate>
<gate>
<ID>656</ID>
<type>FF_GND</type>
<position>516.5,77.5</position>
<output>
<ID>OUT_0</ID>760 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>271</ID>
<type>DE_TO</type>
<position>484,51</position>
<input>
<ID>IN_0</ID>716 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 2</lparam></gate>
<gate>
<ID>273</ID>
<type>DE_TO</type>
<position>486,51</position>
<input>
<ID>IN_0</ID>717 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 3</lparam></gate>
<gate>
<ID>469</ID>
<type>DE_TO</type>
<position>551.5,62</position>
<input>
<ID>IN_0</ID>758 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>277</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>491.5,58</position>
<input>
<ID>ENABLE_0</ID>729 </input>
<input>
<ID>IN_0</ID>580 </input>
<input>
<ID>IN_1</ID>535 </input>
<input>
<ID>IN_2</ID>419 </input>
<input>
<ID>IN_3</ID>578 </input>
<output>
<ID>OUT_0</ID>718 </output>
<output>
<ID>OUT_1</ID>722 </output>
<output>
<ID>OUT_2</ID>723 </output>
<output>
<ID>OUT_3</ID>724 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>279</ID>
<type>DE_TO</type>
<position>489,51</position>
<input>
<ID>IN_0</ID>718 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 4</lparam></gate>
<gate>
<ID>473</ID>
<type>DE_TO</type>
<position>549,61.5</position>
<input>
<ID>IN_0</ID>757 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>474</ID>
<type>DE_TO</type>
<position>546,62</position>
<input>
<ID>IN_0</ID>756 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>481</ID>
<type>DE_TO</type>
<position>542.5,62</position>
<input>
<ID>IN_0</ID>755 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>290</ID>
<type>DE_TO</type>
<position>491,51</position>
<input>
<ID>IN_0</ID>722 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 5</lparam></gate>
<gate>
<ID>484</ID>
<type>DE_TO</type>
<position>540,62</position>
<input>
<ID>IN_0</ID>754 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>292</ID>
<type>DE_TO</type>
<position>493,51</position>
<input>
<ID>IN_0</ID>723 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 6</lparam></gate>
<gate>
<ID>686</ID>
<type>DA_FROM</type>
<position>439,86</position>
<input>
<ID>IN_0</ID>792 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>1074</ID>
<type>AA_LABEL</type>
<position>485.5,108</position>
<gparam>LABEL_TEXT Address Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>688</ID>
<type>DA_FROM</type>
<position>439,83</position>
<input>
<ID>IN_0</ID>793 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>690</ID>
<type>DA_FROM</type>
<position>439,80.5</position>
<input>
<ID>IN_0</ID>794 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>692</ID>
<type>DA_FROM</type>
<position>439,78</position>
<input>
<ID>IN_0</ID>795 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>113</ID>
<type>AI_REGISTER12</type>
<position>476,70</position>
<input>
<ID>IN_0</ID>780 </input>
<input>
<ID>IN_1</ID>775 </input>
<input>
<ID>IN_10</ID>784 </input>
<input>
<ID>IN_11</ID>783 </input>
<input>
<ID>IN_2</ID>776 </input>
<input>
<ID>IN_3</ID>777 </input>
<input>
<ID>IN_4</ID>778 </input>
<input>
<ID>IN_5</ID>779 </input>
<input>
<ID>IN_6</ID>774 </input>
<input>
<ID>IN_7</ID>773 </input>
<input>
<ID>IN_8</ID>782 </input>
<input>
<ID>IN_9</ID>781 </input>
<output>
<ID>OUT_0</ID>622 </output>
<output>
<ID>OUT_1</ID>582 </output>
<output>
<ID>OUT_10</ID>421 </output>
<output>
<ID>OUT_11</ID>420 </output>
<output>
<ID>OUT_2</ID>581 </output>
<output>
<ID>OUT_3</ID>623 </output>
<output>
<ID>OUT_4</ID>580 </output>
<output>
<ID>OUT_5</ID>535 </output>
<output>
<ID>OUT_6</ID>419 </output>
<output>
<ID>OUT_7</ID>578 </output>
<output>
<ID>OUT_8</ID>536 </output>
<output>
<ID>OUT_9</ID>338 </output>
<input>
<ID>clear</ID>300 </input>
<input>
<ID>clock</ID>265 </input>
<input>
<ID>count_enable</ID>337 </input>
<input>
<ID>count_up</ID>305 </input>
<input>
<ID>load</ID>333 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>310</ID>
<type>DE_TO</type>
<position>495,51</position>
<input>
<ID>IN_0</ID>724 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 7</lparam></gate>
<gate>
<ID>311</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>501,58</position>
<input>
<ID>ENABLE_0</ID>729 </input>
<input>
<ID>IN_0</ID>536 </input>
<input>
<ID>IN_1</ID>338 </input>
<input>
<ID>IN_2</ID>421 </input>
<input>
<ID>IN_3</ID>420 </input>
<output>
<ID>OUT_0</ID>725 </output>
<output>
<ID>OUT_1</ID>726 </output>
<output>
<ID>OUT_2</ID>727 </output>
<output>
<ID>OUT_3</ID>728 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>517</ID>
<type>DE_TO</type>
<position>537,62</position>
<input>
<ID>IN_0</ID>753 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>518</ID>
<type>DE_TO</type>
<position>534.5,62</position>
<input>
<ID>IN_0</ID>752 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>520</ID>
<type>DE_TO</type>
<position>512,61.5</position>
<input>
<ID>IN_0</ID>744 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>327</ID>
<type>DE_TO</type>
<position>498.5,51</position>
<input>
<ID>IN_0</ID>725 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 8</lparam></gate>
<gate>
<ID>908</ID>
<type>DA_FROM</type>
<position>574,-10.5</position>
<input>
<ID>IN_0</ID>885 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>909</ID>
<type>DA_FROM</type>
<position>573.5,-13.5</position>
<input>
<ID>IN_0</ID>880 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>910</ID>
<type>DA_FROM</type>
<position>573.5,-16.5</position>
<input>
<ID>IN_0</ID>879 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>911</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>593,-4</position>
<input>
<ID>ENABLE_0</ID>891 </input>
<input>
<ID>IN_0</ID>879 </input>
<input>
<ID>IN_1</ID>880 </input>
<input>
<ID>IN_2</ID>885 </input>
<input>
<ID>IN_3</ID>886 </input>
<input>
<ID>IN_4</ID>887 </input>
<input>
<ID>IN_5</ID>888 </input>
<input>
<ID>IN_6</ID>889 </input>
<input>
<ID>IN_7</ID>890 </input>
<output>
<ID>OUT_0</ID>892 </output>
<output>
<ID>OUT_1</ID>893 </output>
<output>
<ID>OUT_2</ID>894 </output>
<output>
<ID>OUT_3</ID>895 </output>
<output>
<ID>OUT_4</ID>896 </output>
<output>
<ID>OUT_5</ID>897 </output>
<output>
<ID>OUT_6</ID>898 </output>
<output>
<ID>OUT_7</ID>899 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>912</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>588.5,2</position>
<input>
<ID>ENABLE_0</ID>891 </input>
<input>
<ID>IN_0</ID>884 </input>
<input>
<ID>IN_1</ID>883 </input>
<input>
<ID>IN_2</ID>882 </input>
<input>
<ID>IN_3</ID>881 </input>
<output>
<ID>OUT_0</ID>900 </output>
<output>
<ID>OUT_1</ID>901 </output>
<output>
<ID>OUT_2</ID>903 </output>
<output>
<ID>OUT_3</ID>904 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>913</ID>
<type>DA_FROM</type>
<position>574,14</position>
<input>
<ID>IN_0</ID>881 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A11</lparam></gate>
<gate>
<ID>914</ID>
<type>DA_FROM</type>
<position>574,11</position>
<input>
<ID>IN_0</ID>882 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A10</lparam></gate>
<gate>
<ID>915</ID>
<type>DA_FROM</type>
<position>574,8.5</position>
<input>
<ID>IN_0</ID>883 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A9</lparam></gate>
<gate>
<ID>916</ID>
<type>DA_FROM</type>
<position>574,6</position>
<input>
<ID>IN_0</ID>884 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A8</lparam></gate>
<gate>
<ID>530</ID>
<type>DE_TO</type>
<position>515.5,61.5</position>
<input>
<ID>IN_0</ID>745 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>917</ID>
<type>DA_FROM</type>
<position>574,3</position>
<input>
<ID>IN_0</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A7</lparam></gate>
<gate>
<ID>918</ID>
<type>DA_FROM</type>
<position>574,0.5</position>
<input>
<ID>IN_0</ID>889 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A6</lparam></gate>
<gate>
<ID>919</ID>
<type>DA_FROM</type>
<position>574,-2.5</position>
<input>
<ID>IN_0</ID>888 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A5</lparam></gate>
<gate>
<ID>920</ID>
<type>DA_FROM</type>
<position>574,-5</position>
<input>
<ID>IN_0</ID>887 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A4</lparam></gate>
<gate>
<ID>921</ID>
<type>DA_FROM</type>
<position>574,-7.5</position>
<input>
<ID>IN_0</ID>886 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>922</ID>
<type>DE_TO</type>
<position>613.5,-15.5</position>
<input>
<ID>IN_0</ID>892 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Addr 0</lparam></gate>
<gate>
<ID>923</ID>
<type>DE_TO</type>
<position>613,-12.5</position>
<input>
<ID>IN_0</ID>893 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Addr 1</lparam></gate>
<gate>
<ID>151</ID>
<type>DA_FROM</type>
<position>475,57</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>924</ID>
<type>DE_TO</type>
<position>613,-9.5</position>
<input>
<ID>IN_0</ID>894 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Addr 2</lparam></gate>
<gate>
<ID>925</ID>
<type>DE_TO</type>
<position>613,-7</position>
<input>
<ID>IN_0</ID>895 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Addr 3</lparam></gate>
<gate>
<ID>153</ID>
<type>DA_FROM</type>
<position>477,59</position>
<input>
<ID>IN_0</ID>300 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>926</ID>
<type>DE_TO</type>
<position>613,-4.5</position>
<input>
<ID>IN_0</ID>896 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Addr 4</lparam></gate>
<gate>
<ID>927</ID>
<type>DE_TO</type>
<position>613,-2</position>
<input>
<ID>IN_0</ID>897 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Addr 5</lparam></gate>
<gate>
<ID>155</ID>
<type>EE_VDD</type>
<position>477,81</position>
<output>
<ID>OUT_0</ID>305 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>928</ID>
<type>DE_TO</type>
<position>613,0.5</position>
<input>
<ID>IN_0</ID>898 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Addr 6</lparam></gate>
<gate>
<ID>156</ID>
<type>DA_FROM</type>
<position>469,86</position>
<input>
<ID>IN_0</ID>333 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load-ADREG</lparam></gate>
<gate>
<ID>929</ID>
<type>DE_TO</type>
<position>613,3</position>
<input>
<ID>IN_0</ID>899 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Addr 7</lparam></gate>
<gate>
<ID>930</ID>
<type>DE_TO</type>
<position>613,5.5</position>
<input>
<ID>IN_0</ID>900 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Addr 8</lparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>468,89.5</position>
<input>
<ID>IN_0</ID>337 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INC-ADREG</lparam></gate>
<gate>
<ID>931</ID>
<type>DE_TO</type>
<position>613,8</position>
<input>
<ID>IN_0</ID>901 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Addr 9</lparam></gate>
<gate>
<ID>932</ID>
<type>DE_TO</type>
<position>613,10.5</position>
<input>
<ID>IN_0</ID>903 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Addr 10</lparam></gate>
<gate>
<ID>160</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>513.5,72</position>
<input>
<ID>ENABLE_0</ID>628 </input>
<input>
<ID>IN_0</ID>580 </input>
<input>
<ID>IN_1</ID>535 </input>
<input>
<ID>IN_2</ID>419 </input>
<input>
<ID>IN_3</ID>578 </input>
<input>
<ID>IN_4</ID>536 </input>
<input>
<ID>IN_5</ID>338 </input>
<input>
<ID>IN_6</ID>421 </input>
<input>
<ID>IN_7</ID>420 </input>
<output>
<ID>OUT_0</ID>748 </output>
<output>
<ID>OUT_1</ID>749 </output>
<output>
<ID>OUT_2</ID>750 </output>
<output>
<ID>OUT_3</ID>751 </output>
<output>
<ID>OUT_4</ID>752 </output>
<output>
<ID>OUT_5</ID>753 </output>
<output>
<ID>OUT_6</ID>754 </output>
<output>
<ID>OUT_7</ID>755 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>933</ID>
<type>DE_TO</type>
<position>613,13</position>
<input>
<ID>IN_0</ID>904 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Addr 11</lparam></gate>
<gate>
<ID>934</ID>
<type>DA_FROM</type>
<position>590.5,8</position>
<input>
<ID>IN_0</ID>891 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Res-ADDR</lparam></gate>
<gate>
<ID>745</ID>
<type>DA_FROM</type>
<position>439,75</position>
<input>
<ID>IN_0</ID>801 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>363</ID>
<type>DE_TO</type>
<position>500.5,51</position>
<input>
<ID>IN_0</ID>726 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 9</lparam></gate>
<gate>
<ID>751</ID>
<type>DA_FROM</type>
<position>439,72.5</position>
<input>
<ID>IN_0</ID>800 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>367</ID>
<type>DE_TO</type>
<position>502.5,51</position>
<input>
<ID>IN_0</ID>727 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 10</lparam></gate>
<gate>
<ID>754</ID>
<type>DA_FROM</type>
<position>439,69.5</position>
<input>
<ID>IN_0</ID>799 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>756</ID>
<type>DA_FROM</type>
<position>439,67</position>
<input>
<ID>IN_0</ID>798 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>758</ID>
<type>DA_FROM</type>
<position>439,64.5</position>
<input>
<ID>IN_0</ID>797 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>380</ID>
<type>DE_TO</type>
<position>504.5,51</position>
<input>
<ID>IN_0</ID>728 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 11</lparam></gate>
<wire>
<ID>580</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481,68.5,511.5,68.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<connection>
<GID>113</GID>
<name>OUT_4</name></connection>
<intersection>490 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>490,60,490,68.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>68.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>773</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>458.5,71.5,471,71.5</points>
<connection>
<GID>113</GID>
<name>IN_7</name></connection>
<connection>
<GID>798</GID>
<name>OUT_7</name></connection>
<intersection>464 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>464,34.5,464,71.5</points>
<intersection>34.5 7</intersection>
<intersection>71.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>451.5,34.5,464,34.5</points>
<connection>
<GID>815</GID>
<name>OUT_7</name></connection>
<intersection>464 6</intersection></hsegment></shape></wire>
<wire>
<ID>774</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>458.5,70.5,471,70.5</points>
<connection>
<GID>113</GID>
<name>IN_6</name></connection>
<connection>
<GID>798</GID>
<name>OUT_6</name></connection>
<intersection>465 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>465,33.5,465,70.5</points>
<intersection>33.5 7</intersection>
<intersection>70.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>451.5,33.5,465,33.5</points>
<connection>
<GID>815</GID>
<name>OUT_6</name></connection>
<intersection>465 6</intersection></hsegment></shape></wire>
<wire>
<ID>581</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481,66.5,507,66.5</points>
<connection>
<GID>203</GID>
<name>IN_2</name></connection>
<connection>
<GID>113</GID>
<name>OUT_2</name></connection>
<intersection>483 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>483,60,483,66.5</points>
<connection>
<GID>265</GID>
<name>IN_2</name></connection>
<intersection>66.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>775</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>458.5,65.5,471,65.5</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<connection>
<GID>798</GID>
<name>OUT_1</name></connection>
<intersection>470 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>470,28.5,470,65.5</points>
<intersection>28.5 16</intersection>
<intersection>65.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>451.5,28.5,470,28.5</points>
<connection>
<GID>815</GID>
<name>OUT_1</name></connection>
<intersection>470 15</intersection></hsegment></shape></wire>
<wire>
<ID>582</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481,65.5,507,65.5</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<connection>
<GID>113</GID>
<name>OUT_1</name></connection>
<intersection>482 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>482,60,482,65.5</points>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<intersection>65.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>776</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>458.5,66.5,471,66.5</points>
<connection>
<GID>113</GID>
<name>IN_2</name></connection>
<connection>
<GID>798</GID>
<name>OUT_2</name></connection>
<intersection>469 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>469,29.5,469,66.5</points>
<intersection>29.5 16</intersection>
<intersection>66.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>451.5,29.5,469,29.5</points>
<connection>
<GID>815</GID>
<name>OUT_2</name></connection>
<intersection>469 15</intersection></hsegment></shape></wire>
<wire>
<ID>777</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>458.5,67.5,471,67.5</points>
<connection>
<GID>113</GID>
<name>IN_3</name></connection>
<connection>
<GID>798</GID>
<name>OUT_3</name></connection>
<intersection>468 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>468,30.5,468,67.5</points>
<intersection>30.5 16</intersection>
<intersection>67.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>451.5,30.5,468,30.5</points>
<connection>
<GID>815</GID>
<name>OUT_3</name></connection>
<intersection>468 15</intersection></hsegment></shape></wire>
<wire>
<ID>778</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>458.5,68.5,471,68.5</points>
<connection>
<GID>113</GID>
<name>IN_4</name></connection>
<connection>
<GID>798</GID>
<name>OUT_4</name></connection>
<intersection>467 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>467,31.5,467,68.5</points>
<intersection>31.5 10</intersection>
<intersection>68.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>451.5,31.5,467,31.5</points>
<connection>
<GID>815</GID>
<name>OUT_4</name></connection>
<intersection>467 9</intersection></hsegment></shape></wire>
<wire>
<ID>779</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>458.5,69.5,471,69.5</points>
<connection>
<GID>113</GID>
<name>IN_5</name></connection>
<connection>
<GID>798</GID>
<name>OUT_5</name></connection>
<intersection>466 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>466,32.5,466,69.5</points>
<intersection>32.5 10</intersection>
<intersection>69.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>451.5,32.5,466,32.5</points>
<connection>
<GID>815</GID>
<name>OUT_5</name></connection>
<intersection>466 9</intersection></hsegment></shape></wire>
<wire>
<ID>780</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>458.5,64.5,471,64.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<connection>
<GID>798</GID>
<name>OUT_0</name></connection>
<intersection>471 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>471,27.5,471,64.5</points>
<intersection>27.5 16</intersection>
<intersection>64.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>451.5,27.5,471,27.5</points>
<connection>
<GID>815</GID>
<name>OUT_0</name></connection>
<intersection>471 15</intersection></hsegment></shape></wire>
<wire>
<ID>781</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>454.5,73.5,471,73.5</points>
<connection>
<GID>113</GID>
<name>IN_9</name></connection>
<connection>
<GID>800</GID>
<name>OUT_1</name></connection>
<intersection>462 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>462,36.5,462,73.5</points>
<intersection>36.5 7</intersection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>447,36.5,462,36.5</points>
<connection>
<GID>816</GID>
<name>OUT_1</name></connection>
<intersection>462 6</intersection></hsegment></shape></wire>
<wire>
<ID>782</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>454.5,72.5,471,72.5</points>
<connection>
<GID>113</GID>
<name>IN_8</name></connection>
<connection>
<GID>800</GID>
<name>OUT_0</name></connection>
<intersection>463 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>463,35.5,463,72.5</points>
<intersection>35.5 7</intersection>
<intersection>72.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>447,35.5,463,35.5</points>
<connection>
<GID>816</GID>
<name>OUT_0</name></connection>
<intersection>463 6</intersection></hsegment></shape></wire>
<wire>
<ID>783</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>454.5,75.5,471,75.5</points>
<connection>
<GID>113</GID>
<name>IN_11</name></connection>
<connection>
<GID>800</GID>
<name>OUT_3</name></connection>
<intersection>460 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>460,38.5,460,75.5</points>
<intersection>38.5 7</intersection>
<intersection>75.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>447,38.5,460,38.5</points>
<connection>
<GID>816</GID>
<name>OUT_3</name></connection>
<intersection>460 6</intersection></hsegment></shape></wire>
<wire>
<ID>784</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>454.5,74.5,471,74.5</points>
<connection>
<GID>113</GID>
<name>IN_10</name></connection>
<connection>
<GID>800</GID>
<name>OUT_2</name></connection>
<intersection>461 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>461,37.5,461,74.5</points>
<intersection>37.5 7</intersection>
<intersection>74.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>447,37.5,461,37.5</points>
<connection>
<GID>816</GID>
<name>OUT_2</name></connection>
<intersection>461 6</intersection></hsegment></shape></wire>
<wire>
<ID>785</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449,55.5,449,64.5</points>
<intersection>55.5 2</intersection>
<intersection>64.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>440.5,55.5,449,55.5</points>
<connection>
<GID>796</GID>
<name>IN_0</name></connection>
<intersection>449 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>449,64.5,454.5,64.5</points>
<connection>
<GID>798</GID>
<name>IN_0</name></connection>
<intersection>449 0</intersection></hsegment></shape></wire>
<wire>
<ID>786</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448,58.5,448,65.5</points>
<intersection>58.5 2</intersection>
<intersection>65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>448,65.5,454.5,65.5</points>
<connection>
<GID>798</GID>
<name>IN_1</name></connection>
<intersection>448 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>440.5,58.5,448,58.5</points>
<connection>
<GID>795</GID>
<name>IN_0</name></connection>
<intersection>448 0</intersection></hsegment></shape></wire>
<wire>
<ID>792</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>450,75.5,450,86</points>
<intersection>75.5 2</intersection>
<intersection>86 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441,86,450,86</points>
<connection>
<GID>686</GID>
<name>IN_0</name></connection>
<intersection>450 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>450,75.5,450.5,75.5</points>
<connection>
<GID>800</GID>
<name>IN_3</name></connection>
<intersection>450 0</intersection></hsegment></shape></wire>
<wire>
<ID>793</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448.5,74.5,448.5,83</points>
<intersection>74.5 2</intersection>
<intersection>83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441,83,448.5,83</points>
<connection>
<GID>688</GID>
<name>IN_0</name></connection>
<intersection>448.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448.5,74.5,450.5,74.5</points>
<connection>
<GID>800</GID>
<name>IN_2</name></connection>
<intersection>448.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>794</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>447.5,73.5,447.5,80.5</points>
<intersection>73.5 3</intersection>
<intersection>80.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>441,80.5,447.5,80.5</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<intersection>447.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>447.5,73.5,450.5,73.5</points>
<connection>
<GID>800</GID>
<name>IN_1</name></connection>
<intersection>447.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>795</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>446,72.5,446,78</points>
<intersection>72.5 1</intersection>
<intersection>78 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>446,72.5,450.5,72.5</points>
<connection>
<GID>800</GID>
<name>IN_0</name></connection>
<intersection>446 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>441,78,446,78</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<intersection>446 0</intersection></hsegment></shape></wire>
<wire>
<ID>796</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>446.5,61.5,446.5,66.5</points>
<intersection>61.5 3</intersection>
<intersection>66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>446.5,66.5,454.5,66.5</points>
<connection>
<GID>798</GID>
<name>IN_2</name></connection>
<intersection>446.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>441,61.5,446.5,61.5</points>
<connection>
<GID>791</GID>
<name>IN_0</name></connection>
<intersection>446.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>797</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445.5,64.5,445.5,67.5</points>
<intersection>64.5 2</intersection>
<intersection>67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445.5,67.5,454.5,67.5</points>
<connection>
<GID>798</GID>
<name>IN_3</name></connection>
<intersection>445.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>441,64.5,445.5,64.5</points>
<connection>
<GID>758</GID>
<name>IN_0</name></connection>
<intersection>445.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>798</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444,67,444,68.5</points>
<intersection>67 1</intersection>
<intersection>68.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441,67,444,67</points>
<connection>
<GID>756</GID>
<name>IN_0</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444,68.5,454.5,68.5</points>
<connection>
<GID>798</GID>
<name>IN_4</name></connection>
<intersection>444 0</intersection></hsegment></shape></wire>
<wire>
<ID>799</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>441,69.5,454.5,69.5</points>
<connection>
<GID>754</GID>
<name>IN_0</name></connection>
<connection>
<GID>798</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>800</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444,70.5,444,72.5</points>
<intersection>70.5 2</intersection>
<intersection>72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441,72.5,444,72.5</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444,70.5,454.5,70.5</points>
<connection>
<GID>798</GID>
<name>IN_6</name></connection>
<intersection>444 0</intersection></hsegment></shape></wire>
<wire>
<ID>801</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445.5,71.5,445.5,75</points>
<intersection>71.5 2</intersection>
<intersection>75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441,75,445.5,75</points>
<connection>
<GID>745</GID>
<name>IN_0</name></connection>
<intersection>445.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>445.5,71.5,454.5,71.5</points>
<connection>
<GID>798</GID>
<name>IN_7</name></connection>
<intersection>445.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>802</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452.5,77,452.5,80.5</points>
<connection>
<GID>800</GID>
<name>ENABLE_0</name></connection>
<intersection>77 2</intersection>
<intersection>80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>452.5,80.5,455.5,80.5</points>
<connection>
<GID>802</GID>
<name>IN_0</name></connection>
<intersection>452.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>452.5,77,456.5,77</points>
<intersection>452.5 0</intersection>
<intersection>456.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>456.5,73,456.5,77</points>
<connection>
<GID>798</GID>
<name>ENABLE_0</name></connection>
<intersection>77 2</intersection></vsegment></shape></wire>
<wire>
<ID>803</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>440.5,18.5,440.5,27.5</points>
<intersection>18.5 2</intersection>
<intersection>27.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>432,18.5,440.5,18.5</points>
<connection>
<GID>814</GID>
<name>IN_0</name></connection>
<intersection>440.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>440.5,27.5,447.5,27.5</points>
<connection>
<GID>815</GID>
<name>IN_0</name></connection>
<intersection>440.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>804</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>439.5,21.5,439.5,28.5</points>
<intersection>21.5 2</intersection>
<intersection>28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>439.5,28.5,447.5,28.5</points>
<connection>
<GID>815</GID>
<name>IN_1</name></connection>
<intersection>439.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>432,21.5,439.5,21.5</points>
<connection>
<GID>813</GID>
<name>IN_0</name></connection>
<intersection>439.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481,70.5,511.5,70.5</points>
<connection>
<GID>160</GID>
<name>IN_2</name></connection>
<connection>
<GID>113</GID>
<name>OUT_6</name></connection>
<intersection>492 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>492,60,492,70.5</points>
<connection>
<GID>277</GID>
<name>IN_2</name></connection>
<intersection>70.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>805</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>441.5,38.5,441.5,49</points>
<intersection>38.5 2</intersection>
<intersection>49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,49,441.5,49</points>
<connection>
<GID>818</GID>
<name>IN_0</name></connection>
<intersection>441.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>441.5,38.5,443,38.5</points>
<connection>
<GID>816</GID>
<name>IN_3</name></connection>
<intersection>441.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481,75.5,511.5,75.5</points>
<connection>
<GID>160</GID>
<name>IN_7</name></connection>
<connection>
<GID>113</GID>
<name>OUT_11</name></connection>
<intersection>502.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>502.5,60,502.5,75.5</points>
<connection>
<GID>311</GID>
<name>IN_3</name></connection>
<intersection>75.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>806</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>440,37.5,440,46</points>
<intersection>37.5 2</intersection>
<intersection>46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,46,440,46</points>
<connection>
<GID>819</GID>
<name>IN_0</name></connection>
<intersection>440 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>440,37.5,443,37.5</points>
<connection>
<GID>816</GID>
<name>IN_2</name></connection>
<intersection>440 0</intersection></hsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481,74.5,511.5,74.5</points>
<connection>
<GID>160</GID>
<name>IN_6</name></connection>
<connection>
<GID>113</GID>
<name>OUT_10</name></connection>
<intersection>501.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>501.5,60,501.5,74.5</points>
<connection>
<GID>311</GID>
<name>IN_2</name></connection>
<intersection>74.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>807</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>439,36.5,439,43.5</points>
<intersection>36.5 3</intersection>
<intersection>43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>432.5,43.5,439,43.5</points>
<connection>
<GID>820</GID>
<name>IN_0</name></connection>
<intersection>439 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>439,36.5,443,36.5</points>
<connection>
<GID>816</GID>
<name>IN_1</name></connection>
<intersection>439 0</intersection></hsegment></shape></wire>
<wire>
<ID>808</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437.5,35.5,437.5,41</points>
<intersection>35.5 1</intersection>
<intersection>41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>437.5,35.5,443,35.5</points>
<connection>
<GID>816</GID>
<name>IN_0</name></connection>
<intersection>437.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>432.5,41,437.5,41</points>
<connection>
<GID>821</GID>
<name>IN_0</name></connection>
<intersection>437.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>809</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>438,24.5,438,29.5</points>
<intersection>24.5 3</intersection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>438,29.5,447.5,29.5</points>
<connection>
<GID>815</GID>
<name>IN_2</name></connection>
<intersection>438 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>432.5,24.5,438,24.5</points>
<connection>
<GID>811</GID>
<name>IN_0</name></connection>
<intersection>438 0</intersection></hsegment></shape></wire>
<wire>
<ID>810</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437,27.5,437,30.5</points>
<intersection>27.5 2</intersection>
<intersection>30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>437,30.5,447.5,30.5</points>
<connection>
<GID>815</GID>
<name>IN_3</name></connection>
<intersection>437 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>432.5,27.5,437,27.5</points>
<connection>
<GID>827</GID>
<name>IN_0</name></connection>
<intersection>437 0</intersection></hsegment></shape></wire>
<wire>
<ID>811</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>435.5,30,435.5,31.5</points>
<intersection>30 1</intersection>
<intersection>31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,30,435.5,30</points>
<connection>
<GID>826</GID>
<name>IN_0</name></connection>
<intersection>435.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>435.5,31.5,447.5,31.5</points>
<connection>
<GID>815</GID>
<name>IN_4</name></connection>
<intersection>435.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>812</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432.5,32.5,447.5,32.5</points>
<connection>
<GID>825</GID>
<name>IN_0</name></connection>
<connection>
<GID>815</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>813</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>435.5,33.5,435.5,35.5</points>
<intersection>33.5 2</intersection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,35.5,435.5,35.5</points>
<connection>
<GID>824</GID>
<name>IN_0</name></connection>
<intersection>435.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>435.5,33.5,447.5,33.5</points>
<connection>
<GID>815</GID>
<name>IN_6</name></connection>
<intersection>435.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>814</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437,34.5,437,38</points>
<intersection>34.5 2</intersection>
<intersection>38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>432.5,38,437,38</points>
<connection>
<GID>823</GID>
<name>IN_0</name></connection>
<intersection>437 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>437,34.5,447.5,34.5</points>
<connection>
<GID>815</GID>
<name>IN_7</name></connection>
<intersection>437 0</intersection></hsegment></shape></wire>
<wire>
<ID>815</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>445,40,472,40</points>
<connection>
<GID>816</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>817</GID>
<name>IN_0</name></connection>
<intersection>449.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>449.5,36,449.5,40</points>
<connection>
<GID>815</GID>
<name>ENABLE_0</name></connection>
<intersection>40 1</intersection></vsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481,64.5,507,64.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>481 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>481,60,481,64.5</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>64.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481,67.5,507,67.5</points>
<connection>
<GID>203</GID>
<name>IN_3</name></connection>
<connection>
<GID>113</GID>
<name>OUT_3</name></connection>
<intersection>484 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>484,60,484,67.5</points>
<connection>
<GID>265</GID>
<name>IN_3</name></connection>
<intersection>67.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>509,69,509,84</points>
<connection>
<GID>203</GID>
<name>ENABLE_0</name></connection>
<intersection>77 13</intersection>
<intersection>84 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>509,84,519.5,84</points>
<connection>
<GID>655</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>509 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>509,77,513.5,77</points>
<connection>
<GID>160</GID>
<name>ENABLE_0</name></connection>
<intersection>509 0</intersection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>475,59,475,62.5</points>
<connection>
<GID>113</GID>
<name>clock</name></connection>
<connection>
<GID>151</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>879</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>584,-16.5,584,-7.5</points>
<intersection>-16.5 2</intersection>
<intersection>-7.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>575.5,-16.5,584,-16.5</points>
<connection>
<GID>910</GID>
<name>IN_0</name></connection>
<intersection>584 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>584,-7.5,591,-7.5</points>
<connection>
<GID>911</GID>
<name>IN_0</name></connection>
<intersection>584 0</intersection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>477,61,477,62.5</points>
<connection>
<GID>113</GID>
<name>clear</name></connection>
<connection>
<GID>153</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>880</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583,-13.5,583,-6.5</points>
<intersection>-13.5 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>583,-6.5,591,-6.5</points>
<connection>
<GID>911</GID>
<name>IN_1</name></connection>
<intersection>583 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>575.5,-13.5,583,-13.5</points>
<connection>
<GID>909</GID>
<name>IN_0</name></connection>
<intersection>583 0</intersection></hsegment></shape></wire>
<wire>
<ID>881</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585,3.5,585,14</points>
<intersection>3.5 2</intersection>
<intersection>14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>576,14,585,14</points>
<connection>
<GID>913</GID>
<name>IN_0</name></connection>
<intersection>585 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>585,3.5,586.5,3.5</points>
<connection>
<GID>912</GID>
<name>IN_3</name></connection>
<intersection>585 0</intersection></hsegment></shape></wire>
<wire>
<ID>882</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583.5,2.5,583.5,11</points>
<intersection>2.5 2</intersection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>576,11,583.5,11</points>
<connection>
<GID>914</GID>
<name>IN_0</name></connection>
<intersection>583.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>583.5,2.5,586.5,2.5</points>
<connection>
<GID>912</GID>
<name>IN_2</name></connection>
<intersection>583.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>883</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>582.5,1.5,582.5,8.5</points>
<intersection>1.5 3</intersection>
<intersection>8.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>576,8.5,582.5,8.5</points>
<connection>
<GID>915</GID>
<name>IN_0</name></connection>
<intersection>582.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>582.5,1.5,586.5,1.5</points>
<connection>
<GID>912</GID>
<name>IN_1</name></connection>
<intersection>582.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>884</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>581,0.5,581,6</points>
<intersection>0.5 1</intersection>
<intersection>6 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>581,0.5,586.5,0.5</points>
<connection>
<GID>912</GID>
<name>IN_0</name></connection>
<intersection>581 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>576,6,581,6</points>
<connection>
<GID>916</GID>
<name>IN_0</name></connection>
<intersection>581 0</intersection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>477,77.5,477,80</points>
<connection>
<GID>113</GID>
<name>count_up</name></connection>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>885</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>581.5,-10.5,581.5,-5.5</points>
<intersection>-10.5 3</intersection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>581.5,-5.5,591,-5.5</points>
<connection>
<GID>911</GID>
<name>IN_2</name></connection>
<intersection>581.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>576,-10.5,581.5,-10.5</points>
<connection>
<GID>908</GID>
<name>IN_0</name></connection>
<intersection>581.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>886</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>580.5,-7.5,580.5,-4.5</points>
<intersection>-7.5 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>580.5,-4.5,591,-4.5</points>
<connection>
<GID>911</GID>
<name>IN_3</name></connection>
<intersection>580.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>576,-7.5,580.5,-7.5</points>
<connection>
<GID>921</GID>
<name>IN_0</name></connection>
<intersection>580.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>887</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>579,-5,579,-3.5</points>
<intersection>-5 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>576,-5,579,-5</points>
<connection>
<GID>920</GID>
<name>IN_0</name></connection>
<intersection>579 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>579,-3.5,591,-3.5</points>
<connection>
<GID>911</GID>
<name>IN_4</name></connection>
<intersection>579 0</intersection></hsegment></shape></wire>
<wire>
<ID>888</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>576,-2.5,591,-2.5</points>
<connection>
<GID>911</GID>
<name>IN_5</name></connection>
<connection>
<GID>919</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>889</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>579,-1.5,579,0.5</points>
<intersection>-1.5 2</intersection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>576,0.5,579,0.5</points>
<connection>
<GID>918</GID>
<name>IN_0</name></connection>
<intersection>579 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>579,-1.5,591,-1.5</points>
<connection>
<GID>911</GID>
<name>IN_6</name></connection>
<intersection>579 0</intersection></hsegment></shape></wire>
<wire>
<ID>890</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>580.5,-0.5,580.5,3</points>
<intersection>-0.5 2</intersection>
<intersection>3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>576,3,580.5,3</points>
<connection>
<GID>917</GID>
<name>IN_0</name></connection>
<intersection>580.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>580.5,-0.5,591,-0.5</points>
<connection>
<GID>911</GID>
<name>IN_7</name></connection>
<intersection>580.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>891</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>588.5,5,593,5</points>
<connection>
<GID>912</GID>
<name>ENABLE_0</name></connection>
<intersection>590.5 5</intersection>
<intersection>593 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>593,1,593,5</points>
<connection>
<GID>911</GID>
<name>ENABLE_0</name></connection>
<intersection>5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>590.5,5,590.5,6</points>
<connection>
<GID>934</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment></shape></wire>
<wire>
<ID>892</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>596.5,-15.5,596.5,-7.5</points>
<intersection>-15.5 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>596.5,-15.5,611.5,-15.5</points>
<connection>
<GID>922</GID>
<name>IN_0</name></connection>
<intersection>596.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>595,-7.5,596.5,-7.5</points>
<connection>
<GID>911</GID>
<name>OUT_0</name></connection>
<intersection>596.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>893</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>597.5,-12.5,597.5,-6.5</points>
<intersection>-12.5 1</intersection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>597.5,-12.5,611,-12.5</points>
<connection>
<GID>923</GID>
<name>IN_0</name></connection>
<intersection>597.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>595,-6.5,597.5,-6.5</points>
<connection>
<GID>911</GID>
<name>OUT_1</name></connection>
<intersection>597.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>894</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>598,-9.5,598,-5.5</points>
<intersection>-9.5 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>598,-9.5,611,-9.5</points>
<connection>
<GID>924</GID>
<name>IN_0</name></connection>
<intersection>598 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>595,-5.5,598,-5.5</points>
<connection>
<GID>911</GID>
<name>OUT_2</name></connection>
<intersection>598 0</intersection></hsegment></shape></wire>
<wire>
<ID>895</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>599.5,-7,599.5,-4.5</points>
<intersection>-7 1</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>599.5,-7,611,-7</points>
<connection>
<GID>925</GID>
<name>IN_0</name></connection>
<intersection>599.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>595,-4.5,599.5,-4.5</points>
<connection>
<GID>911</GID>
<name>OUT_3</name></connection>
<intersection>599.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>896</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>603,-4.5,603,-3.5</points>
<intersection>-4.5 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>603,-4.5,611,-4.5</points>
<connection>
<GID>926</GID>
<name>IN_0</name></connection>
<intersection>603 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>595,-3.5,603,-3.5</points>
<connection>
<GID>911</GID>
<name>OUT_4</name></connection>
<intersection>603 0</intersection></hsegment></shape></wire>
<wire>
<ID>897</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>603,-2.5,603,-2</points>
<intersection>-2.5 1</intersection>
<intersection>-2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>595,-2.5,603,-2.5</points>
<connection>
<GID>911</GID>
<name>OUT_5</name></connection>
<intersection>603 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>603,-2,611,-2</points>
<connection>
<GID>927</GID>
<name>IN_0</name></connection>
<intersection>603 0</intersection></hsegment></shape></wire>
<wire>
<ID>898</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>607,-1.5,607,0.5</points>
<intersection>-1.5 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>595,-1.5,607,-1.5</points>
<connection>
<GID>911</GID>
<name>OUT_6</name></connection>
<intersection>607 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>607,0.5,611,0.5</points>
<connection>
<GID>928</GID>
<name>IN_0</name></connection>
<intersection>607 0</intersection></hsegment></shape></wire>
<wire>
<ID>899</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>606.5,-0.5,606.5,3</points>
<intersection>-0.5 1</intersection>
<intersection>3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>595,-0.5,606.5,-0.5</points>
<connection>
<GID>911</GID>
<name>OUT_7</name></connection>
<intersection>606.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>606.5,3,611,3</points>
<connection>
<GID>929</GID>
<name>IN_0</name></connection>
<intersection>606.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>900</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>600.5,0.5,600.5,5.5</points>
<intersection>0.5 2</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>600.5,5.5,611,5.5</points>
<connection>
<GID>930</GID>
<name>IN_0</name></connection>
<intersection>600.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>590.5,0.5,600.5,0.5</points>
<connection>
<GID>912</GID>
<name>OUT_0</name></connection>
<intersection>600.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>901</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>598,1.5,598,8</points>
<intersection>1.5 2</intersection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>598,8,611,8</points>
<connection>
<GID>931</GID>
<name>IN_0</name></connection>
<intersection>598 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>590.5,1.5,598,1.5</points>
<connection>
<GID>912</GID>
<name>OUT_1</name></connection>
<intersection>598 0</intersection></hsegment></shape></wire>
<wire>
<ID>903</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>597,2.5,597,10.5</points>
<intersection>2.5 2</intersection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>597,10.5,611,10.5</points>
<connection>
<GID>932</GID>
<name>IN_0</name></connection>
<intersection>597 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>590.5,2.5,597,2.5</points>
<connection>
<GID>912</GID>
<name>OUT_2</name></connection>
<intersection>597 0</intersection></hsegment></shape></wire>
<wire>
<ID>904</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>596,3.5,596,13</points>
<intersection>3.5 2</intersection>
<intersection>13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>596,13,611,13</points>
<connection>
<GID>933</GID>
<name>IN_0</name></connection>
<intersection>596 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>590.5,3.5,596,3.5</points>
<connection>
<GID>912</GID>
<name>OUT_3</name></connection>
<intersection>596 0</intersection></hsegment></shape></wire>
<wire>
<ID>714</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>479.5,53,479.5,56</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>56 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>479.5,56,481,56</points>
<connection>
<GID>265</GID>
<name>OUT_0</name></connection>
<intersection>479.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>715</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>482,53,482,56</points>
<connection>
<GID>265</GID>
<name>OUT_1</name></connection>
<connection>
<GID>269</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>716</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484,53,484,56</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>56 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>483,56,484,56</points>
<connection>
<GID>265</GID>
<name>OUT_2</name></connection>
<intersection>484 0</intersection></hsegment></shape></wire>
<wire>
<ID>717</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484,55.5,484,56</points>
<connection>
<GID>265</GID>
<name>OUT_3</name></connection>
<intersection>55.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>486,53,486,55.5</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>55.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>484,55.5,486,55.5</points>
<intersection>484 0</intersection>
<intersection>486 1</intersection></hsegment></shape></wire>
<wire>
<ID>718</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>489,53,489,56</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>56 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>489,56,490,56</points>
<connection>
<GID>277</GID>
<name>OUT_0</name></connection>
<intersection>489 0</intersection></hsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>475,77.5,475,86</points>
<connection>
<GID>113</GID>
<name>load</name></connection>
<intersection>86 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>471,86,475,86</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>475 0</intersection></hsegment></shape></wire>
<wire>
<ID>722</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491,53,491,56</points>
<connection>
<GID>277</GID>
<name>OUT_1</name></connection>
<connection>
<GID>290</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>476,77.5,476,89.5</points>
<connection>
<GID>113</GID>
<name>count_enable</name></connection>
<intersection>89.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>470,89.5,476,89.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>476 0</intersection></hsegment></shape></wire>
<wire>
<ID>723</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>493,53,493,54.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>54.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>492,54.5,493,54.5</points>
<intersection>492 5</intersection>
<intersection>493 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>492,54.5,492,56</points>
<connection>
<GID>277</GID>
<name>OUT_2</name></connection>
<intersection>54.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481,73.5,511.5,73.5</points>
<connection>
<GID>160</GID>
<name>IN_5</name></connection>
<connection>
<GID>113</GID>
<name>OUT_9</name></connection>
<intersection>500.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>500.5,60,500.5,73.5</points>
<connection>
<GID>311</GID>
<name>IN_1</name></connection>
<intersection>73.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>724</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>495,53,495,56</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>56 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>493,56,495,56</points>
<connection>
<GID>277</GID>
<name>OUT_3</name></connection>
<intersection>495 1</intersection></hsegment></shape></wire>
<wire>
<ID>725</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>498.5,53,498.5,56</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>56 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>498.5,56,499.5,56</points>
<connection>
<GID>311</GID>
<name>OUT_0</name></connection>
<intersection>498.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>726</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>500.5,53,500.5,56</points>
<connection>
<GID>311</GID>
<name>OUT_1</name></connection>
<connection>
<GID>363</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>727</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502.5,53,502.5,56</points>
<connection>
<GID>367</GID>
<name>IN_0</name></connection>
<intersection>56 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>501.5,56,502.5,56</points>
<connection>
<GID>311</GID>
<name>OUT_2</name></connection>
<intersection>502.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>728</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502.5,55.5,502.5,56</points>
<connection>
<GID>311</GID>
<name>OUT_3</name></connection>
<intersection>55.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>504.5,53,504.5,55.5</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>55.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>502.5,55.5,504.5,55.5</points>
<intersection>502.5 0</intersection>
<intersection>504.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481,69.5,511.5,69.5</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<connection>
<GID>113</GID>
<name>OUT_5</name></connection>
<intersection>491 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>491,60,491,69.5</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>69.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481,72.5,511.5,72.5</points>
<connection>
<GID>160</GID>
<name>IN_4</name></connection>
<connection>
<GID>113</GID>
<name>OUT_8</name></connection>
<intersection>499.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>499.5,60,499.5,72.5</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>72.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>729</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>509,50.5,510,50.5</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>509 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>509,50.5,509,58</points>
<intersection>50.5 1</intersection>
<intersection>58 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>485.5,58,509,58</points>
<connection>
<GID>265</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>277</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>311</GID>
<name>ENABLE_0</name></connection>
<intersection>509 8</intersection></hsegment></shape></wire>
<wire>
<ID>744</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>511,64.5,512,64.5</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<intersection>512 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>512,63.5,512,64.5</points>
<connection>
<GID>520</GID>
<name>IN_0</name></connection>
<intersection>64.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>745</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>515.5,63.5,515.5,65.5</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<intersection>65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,65.5,515.5,65.5</points>
<connection>
<GID>203</GID>
<name>OUT_1</name></connection>
<intersection>515.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>746</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>518.5,63.5,518.5,66.5</points>
<connection>
<GID>607</GID>
<name>IN_0</name></connection>
<intersection>66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,66.5,518.5,66.5</points>
<connection>
<GID>203</GID>
<name>OUT_2</name></connection>
<intersection>518.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>747</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>521.5,63.5,521.5,67.5</points>
<connection>
<GID>609</GID>
<name>IN_0</name></connection>
<intersection>67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,67.5,521.5,67.5</points>
<connection>
<GID>203</GID>
<name>OUT_3</name></connection>
<intersection>521.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>748</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>524.5,63.5,524.5,68.5</points>
<connection>
<GID>620</GID>
<name>IN_0</name></connection>
<intersection>68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515.5,68.5,524.5,68.5</points>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection>
<intersection>524.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>749</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>527,63.5,527,69.5</points>
<connection>
<GID>632</GID>
<name>IN_0</name></connection>
<intersection>69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515.5,69.5,527,69.5</points>
<connection>
<GID>160</GID>
<name>OUT_1</name></connection>
<intersection>527 0</intersection></hsegment></shape></wire>
<wire>
<ID>750</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>529.5,64,529.5,70.5</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515.5,70.5,529.5,70.5</points>
<connection>
<GID>160</GID>
<name>OUT_2</name></connection>
<intersection>529.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>751</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>531.5,64,531.5,71.5</points>
<connection>
<GID>654</GID>
<name>IN_0</name></connection>
<intersection>71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515.5,71.5,531.5,71.5</points>
<connection>
<GID>160</GID>
<name>OUT_3</name></connection>
<intersection>531.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>752</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>534.5,64,534.5,72.5</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<intersection>72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515.5,72.5,534.5,72.5</points>
<connection>
<GID>160</GID>
<name>OUT_4</name></connection>
<intersection>534.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>753</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>537,64,537,73.5</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515.5,73.5,537,73.5</points>
<connection>
<GID>160</GID>
<name>OUT_5</name></connection>
<intersection>537 0</intersection></hsegment></shape></wire>
<wire>
<ID>754</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540,64,540,74.5</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<intersection>74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515.5,74.5,540,74.5</points>
<connection>
<GID>160</GID>
<name>OUT_6</name></connection>
<intersection>540 0</intersection></hsegment></shape></wire>
<wire>
<ID>755</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>542.5,64,542.5,75.5</points>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<intersection>75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515.5,75.5,542.5,75.5</points>
<connection>
<GID>160</GID>
<name>OUT_7</name></connection>
<intersection>542.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>756</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,64,546,79.5</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<intersection>79.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>521.5,79.5,546,79.5</points>
<connection>
<GID>655</GID>
<name>OUT_0</name></connection>
<intersection>546 0</intersection></hsegment></shape></wire>
<wire>
<ID>757</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>549,63.5,549,80.5</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<intersection>80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>521.5,80.5,549,80.5</points>
<connection>
<GID>655</GID>
<name>OUT_1</name></connection>
<intersection>549 0</intersection></hsegment></shape></wire>
<wire>
<ID>758</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>551.5,64,551.5,81.5</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>81.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>521.5,81.5,551.5,81.5</points>
<connection>
<GID>655</GID>
<name>OUT_2</name></connection>
<intersection>551.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>759</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>554.5,63.5,554.5,82.5</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<intersection>82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>521.5,82.5,554.5,82.5</points>
<connection>
<GID>655</GID>
<name>OUT_3</name></connection>
<intersection>554.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>760</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516.5,78.5,516.5,79.5</points>
<connection>
<GID>656</GID>
<name>OUT_0</name></connection>
<intersection>79.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>516.5,79.5,517.5,79.5</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<intersection>516.5 0</intersection>
<intersection>517.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>517.5,79.5,517.5,82.5</points>
<connection>
<GID>655</GID>
<name>IN_3</name></connection>
<connection>
<GID>655</GID>
<name>IN_2</name></connection>
<connection>
<GID>655</GID>
<name>IN_1</name></connection>
<intersection>79.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>578</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481,71.5,511.5,71.5</points>
<connection>
<GID>160</GID>
<name>IN_3</name></connection>
<connection>
<GID>113</GID>
<name>OUT_7</name></connection>
<intersection>493 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>493,60,493,71.5</points>
<connection>
<GID>277</GID>
<name>IN_3</name></connection>
<intersection>71.5 1</intersection></vsegment></shape></wire></page 6>
<page 7>
<PageViewport>360.411,525.616,1486.41,-120.384</PageViewport>
<gate>
<ID>965</ID>
<type>DE_TO</type>
<position>494,309</position>
<input>
<ID>IN_0</ID>918 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>1</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>491,313.5</position>
<input>
<ID>ENABLE_0</ID>870 </input>
<input>
<ID>IN_0</ID>790 </input>
<input>
<ID>IN_1</ID>789 </input>
<input>
<ID>IN_2</ID>788 </input>
<input>
<ID>IN_3</ID>791 </input>
<output>
<ID>OUT_0</ID>918 </output>
<output>
<ID>OUT_1</ID>919 </output>
<output>
<ID>OUT_2</ID>920 </output>
<output>
<ID>OUT_3</ID>921 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>966</ID>
<type>DE_TO</type>
<position>497.5,309</position>
<input>
<ID>IN_0</ID>919 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>967</ID>
<type>DA_FROM</type>
<position>457,306</position>
<input>
<ID>IN_0</ID>761 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>968</ID>
<type>DA_FROM</type>
<position>459,306.5</position>
<input>
<ID>IN_0</ID>762 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>970</ID>
<type>DA_FROM</type>
<position>451,333.5</position>
<input>
<ID>IN_0</ID>764 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load-SP</lparam></gate>
<gate>
<ID>971</ID>
<type>DA_FROM</type>
<position>450,337</position>
<input>
<ID>IN_0</ID>765 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INC-SP</lparam></gate>
<gate>
<ID>972</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>495.5,319.5</position>
<input>
<ID>ENABLE_0</ID>870 </input>
<input>
<ID>IN_0</ID>787 </input>
<input>
<ID>IN_1</ID>770 </input>
<input>
<ID>IN_2</ID>767 </input>
<input>
<ID>IN_3</ID>772 </input>
<input>
<ID>IN_4</ID>771 </input>
<input>
<ID>IN_5</ID>766 </input>
<input>
<ID>IN_6</ID>769 </input>
<input>
<ID>IN_7</ID>768 </input>
<output>
<ID>OUT_0</ID>922 </output>
<output>
<ID>OUT_1</ID>923 </output>
<output>
<ID>OUT_2</ID>924 </output>
<output>
<ID>OUT_3</ID>925 </output>
<output>
<ID>OUT_4</ID>926 </output>
<output>
<ID>OUT_5</ID>927 </output>
<output>
<ID>OUT_6</ID>928 </output>
<output>
<ID>OUT_7</ID>929 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>973</ID>
<type>DA_FROM</type>
<position>421,322.5</position>
<input>
<ID>IN_0</ID>958 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>974</ID>
<type>DE_TO</type>
<position>471.5,278.5</position>
<input>
<ID>IN_0</ID>995 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 9</lparam></gate>
<gate>
<ID>10</ID>
<type>DA_FROM</type>
<position>421,309</position>
<input>
<ID>IN_0</ID>953 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>975</ID>
<type>DA_FROM</type>
<position>421,320</position>
<input>
<ID>IN_0</ID>957 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>976</ID>
<type>DE_TO</type>
<position>468,278.5</position>
<input>
<ID>IN_0</ID>994 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 10</lparam></gate>
<gate>
<ID>977</ID>
<type>DA_FROM</type>
<position>421,317</position>
<input>
<ID>IN_0</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>978</ID>
<type>DA_FROM</type>
<position>421,314.5</position>
<input>
<ID>IN_0</ID>955 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>979</ID>
<type>DA_FROM</type>
<position>421,312</position>
<input>
<ID>IN_0</ID>954 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>980</ID>
<type>DE_TO</type>
<position>465,278.5</position>
<input>
<ID>IN_0</ID>993 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 11</lparam></gate>
<gate>
<ID>984</ID>
<type>AE_FULLADDER_4BIT</type>
<position>468.5,292</position>
<input>
<ID>IN_0</ID>771 </input>
<input>
<ID>IN_1</ID>766 </input>
<input>
<ID>IN_2</ID>769 </input>
<input>
<ID>IN_3</ID>768 </input>
<input>
<ID>IN_B_0</ID>1001 </input>
<input>
<ID>IN_B_1</ID>1001 </input>
<input>
<ID>IN_B_2</ID>1001 </input>
<input>
<ID>IN_B_3</ID>1001 </input>
<output>
<ID>OUT_0</ID>984 </output>
<output>
<ID>OUT_1</ID>986 </output>
<output>
<ID>OUT_2</ID>987 </output>
<output>
<ID>OUT_3</ID>985 </output>
<input>
<ID>carry_in</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>986</ID>
<type>AE_FULLADDER_4BIT</type>
<position>485,292</position>
<input>
<ID>IN_0</ID>787 </input>
<input>
<ID>IN_1</ID>770 </input>
<input>
<ID>IN_2</ID>767 </input>
<input>
<ID>IN_3</ID>772 </input>
<input>
<ID>IN_B_0</ID>1001 </input>
<input>
<ID>IN_B_1</ID>1001 </input>
<input>
<ID>IN_B_2</ID>1001 </input>
<input>
<ID>IN_B_3</ID>1001 </input>
<output>
<ID>OUT_0</ID>982 </output>
<output>
<ID>OUT_1</ID>983 </output>
<output>
<ID>OUT_2</ID>981 </output>
<output>
<ID>OUT_3</ID>980 </output>
<input>
<ID>carry_in</ID>973 </input>
<output>
<ID>carry_out</ID>974 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>988</ID>
<type>AE_FULLADDER_4BIT</type>
<position>501.5,292</position>
<input>
<ID>IN_0</ID>790 </input>
<input>
<ID>IN_1</ID>789 </input>
<input>
<ID>IN_2</ID>788 </input>
<input>
<ID>IN_3</ID>791 </input>
<input>
<ID>IN_B_0</ID>1001 </input>
<input>
<ID>IN_B_1</ID>1001 </input>
<input>
<ID>IN_B_2</ID>1001 </input>
<input>
<ID>IN_B_3</ID>1001 </input>
<output>
<ID>OUT_0</ID>976 </output>
<output>
<ID>OUT_1</ID>977 </output>
<output>
<ID>OUT_2</ID>978 </output>
<output>
<ID>OUT_3</ID>979 </output>
<input>
<ID>carry_in</ID>975 </input>
<output>
<ID>carry_out</ID>973 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>797</ID>
<type>DA_FROM</type>
<position>412,266</position>
<input>
<ID>IN_0</ID>960 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>990</ID>
<type>FF_GND</type>
<position>510.5,291</position>
<output>
<ID>OUT_0</ID>975 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>799</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>431.5,278.5</position>
<input>
<ID>ENABLE_0</ID>972 </input>
<input>
<ID>IN_0</ID>960 </input>
<input>
<ID>IN_1</ID>961 </input>
<input>
<ID>IN_2</ID>966 </input>
<input>
<ID>IN_3</ID>967 </input>
<input>
<ID>IN_4</ID>968 </input>
<input>
<ID>IN_5</ID>969 </input>
<input>
<ID>IN_6</ID>970 </input>
<input>
<ID>IN_7</ID>971 </input>
<output>
<ID>OUT_0</ID>942 </output>
<output>
<ID>OUT_1</ID>937 </output>
<output>
<ID>OUT_2</ID>938 </output>
<output>
<ID>OUT_3</ID>939 </output>
<output>
<ID>OUT_4</ID>940 </output>
<output>
<ID>OUT_5</ID>941 </output>
<output>
<ID>OUT_6</ID>936 </output>
<output>
<ID>OUT_7</ID>935 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>992</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>501.5,285</position>
<input>
<ID>ENABLE_0</ID>988 </input>
<input>
<ID>IN_0</ID>979 </input>
<input>
<ID>IN_1</ID>978 </input>
<input>
<ID>IN_2</ID>977 </input>
<input>
<ID>IN_3</ID>976 </input>
<output>
<ID>OUT_0</ID>992 </output>
<output>
<ID>OUT_1</ID>991 </output>
<output>
<ID>OUT_2</ID>990 </output>
<output>
<ID>OUT_3</ID>989 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>801</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>427,284.5</position>
<input>
<ID>ENABLE_0</ID>972 </input>
<input>
<ID>IN_0</ID>965 </input>
<input>
<ID>IN_1</ID>964 </input>
<input>
<ID>IN_2</ID>963 </input>
<input>
<ID>IN_3</ID>962 </input>
<output>
<ID>OUT_0</ID>944 </output>
<output>
<ID>OUT_1</ID>943 </output>
<output>
<ID>OUT_2</ID>946 </output>
<output>
<ID>OUT_3</ID>945 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>994</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>485,285</position>
<input>
<ID>ENABLE_0</ID>988 </input>
<input>
<ID>IN_0</ID>980 </input>
<input>
<ID>IN_1</ID>981 </input>
<input>
<ID>IN_2</ID>983 </input>
<input>
<ID>IN_3</ID>982 </input>
<output>
<ID>OUT_0</ID>1000 </output>
<output>
<ID>OUT_1</ID>999 </output>
<output>
<ID>OUT_2</ID>998 </output>
<output>
<ID>OUT_3</ID>997 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>996</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>468.5,285</position>
<input>
<ID>ENABLE_0</ID>988 </input>
<input>
<ID>IN_0</ID>985 </input>
<input>
<ID>IN_1</ID>987 </input>
<input>
<ID>IN_2</ID>986 </input>
<input>
<ID>IN_3</ID>984 </input>
<output>
<ID>OUT_0</ID>993 </output>
<output>
<ID>OUT_1</ID>994 </output>
<output>
<ID>OUT_2</ID>995 </output>
<output>
<ID>OUT_3</ID>996 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>998</ID>
<type>DA_FROM</type>
<position>516,296.5</position>
<input>
<ID>IN_0</ID>1001 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SP-DEC</lparam></gate>
<gate>
<ID>999</ID>
<type>DA_FROM</type>
<position>471.5,327.5</position>
<input>
<ID>IN_0</ID>1002 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SP-DEC</lparam></gate>
<gate>
<ID>1001</ID>
<type>AE_SMALL_INVERTER</type>
<position>467.5,327.5</position>
<input>
<ID>IN_0</ID>1002 </input>
<output>
<ID>OUT_0</ID>1003 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>822</ID>
<type>DA_FROM</type>
<position>433,289.5</position>
<input>
<ID>IN_0</ID>972 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID RES-SP</lparam></gate>
<gate>
<ID>828</ID>
<type>DA_FROM</type>
<position>412.5,296.5</position>
<input>
<ID>IN_0</ID>962 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A11</lparam></gate>
<gate>
<ID>657</ID>
<type>DA_FROM</type>
<position>420.5,306</position>
<input>
<ID>IN_0</ID>948 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>658</ID>
<type>DA_FROM</type>
<position>420.5,303</position>
<input>
<ID>IN_0</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>659</ID>
<type>DA_FROM</type>
<position>510,285</position>
<input>
<ID>IN_0</ID>988 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SP-ADDR</lparam></gate>
<gate>
<ID>661</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>438.5,315.5</position>
<input>
<ID>ENABLE_0</ID>959 </input>
<input>
<ID>IN_0</ID>947 </input>
<input>
<ID>IN_1</ID>948 </input>
<input>
<ID>IN_2</ID>953 </input>
<input>
<ID>IN_3</ID>954 </input>
<input>
<ID>IN_4</ID>955 </input>
<input>
<ID>IN_5</ID>956 </input>
<input>
<ID>IN_6</ID>957 </input>
<input>
<ID>IN_7</ID>958 </input>
<output>
<ID>OUT_0</ID>942 </output>
<output>
<ID>OUT_1</ID>937 </output>
<output>
<ID>OUT_2</ID>938 </output>
<output>
<ID>OUT_3</ID>939 </output>
<output>
<ID>OUT_4</ID>940 </output>
<output>
<ID>OUT_5</ID>941 </output>
<output>
<ID>OUT_6</ID>936 </output>
<output>
<ID>OUT_7</ID>935 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>663</ID>
<type>DE_TO</type>
<position>536.5,309</position>
<input>
<ID>IN_0</ID>933 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>665</ID>
<type>DE_TO</type>
<position>500.5,309</position>
<input>
<ID>IN_0</ID>920 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>667</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>434.5,321.5</position>
<input>
<ID>ENABLE_0</ID>959 </input>
<input>
<ID>IN_0</ID>952 </input>
<input>
<ID>IN_1</ID>951 </input>
<input>
<ID>IN_2</ID>950 </input>
<input>
<ID>IN_3</ID>949 </input>
<output>
<ID>OUT_0</ID>944 </output>
<output>
<ID>OUT_1</ID>943 </output>
<output>
<ID>OUT_2</ID>946 </output>
<output>
<ID>OUT_3</ID>945 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>676</ID>
<type>DE_TO</type>
<position>503.5,309</position>
<input>
<ID>IN_0</ID>921 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>870</ID>
<type>DA_FROM</type>
<position>412.5,293.5</position>
<input>
<ID>IN_0</ID>963 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A10</lparam></gate>
<gate>
<ID>678</ID>
<type>DA_FROM</type>
<position>439.5,328</position>
<input>
<ID>IN_0</ID>959 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID BUS-SP</lparam></gate>
<gate>
<ID>871</ID>
<type>DA_FROM</type>
<position>412.5,291</position>
<input>
<ID>IN_0</ID>964 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A9</lparam></gate>
<gate>
<ID>872</ID>
<type>DA_FROM</type>
<position>412.5,288.5</position>
<input>
<ID>IN_0</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A8</lparam></gate>
<gate>
<ID>680</ID>
<type>DA_FROM</type>
<position>412.5,272</position>
<input>
<ID>IN_0</ID>966 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>873</ID>
<type>DA_FROM</type>
<position>412.5,285.5</position>
<input>
<ID>IN_0</ID>971 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A7</lparam></gate>
<gate>
<ID>874</ID>
<type>DA_FROM</type>
<position>412.5,283</position>
<input>
<ID>IN_0</ID>970 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A6</lparam></gate>
<gate>
<ID>682</ID>
<type>DE_TO</type>
<position>506.5,309</position>
<input>
<ID>IN_0</ID>922 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>684</ID>
<type>DA_FROM</type>
<position>412,269</position>
<input>
<ID>IN_0</ID>961 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>885</ID>
<type>DE_TO</type>
<position>509,309</position>
<input>
<ID>IN_0</ID>923 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>896</ID>
<type>DA_FROM</type>
<position>412.5,280</position>
<input>
<ID>IN_0</ID>969 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A5</lparam></gate>
<gate>
<ID>897</ID>
<type>DA_FROM</type>
<position>412.5,277.5</position>
<input>
<ID>IN_0</ID>968 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A4</lparam></gate>
<gate>
<ID>898</ID>
<type>DA_FROM</type>
<position>412.5,275</position>
<input>
<ID>IN_0</ID>967 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>899</ID>
<type>DA_FROM</type>
<position>489,331.5</position>
<input>
<ID>IN_0</ID>870 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SP-BUS</lparam></gate>
<gate>
<ID>901</ID>
<type>DE_TO</type>
<position>505,278.5</position>
<input>
<ID>IN_0</ID>989 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 0</lparam></gate>
<gate>
<ID>902</ID>
<type>DE_TO</type>
<position>511.5,309.5</position>
<input>
<ID>IN_0</ID>924 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>903</ID>
<type>DE_TO</type>
<position>513.5,309.5</position>
<input>
<ID>IN_0</ID>925 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>904</ID>
<type>DE_TO</type>
<position>502,278</position>
<input>
<ID>IN_0</ID>990 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 1</lparam></gate>
<gate>
<ID>905</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>501.5,328.5</position>
<input>
<ID>ENABLE_0</ID>870 </input>
<input>
<ID>IN_0</ID>934 </input>
<input>
<ID>IN_1</ID>934 </input>
<input>
<ID>IN_2</ID>934 </input>
<input>
<ID>IN_3</ID>934 </input>
<output>
<ID>OUT_0</ID>930 </output>
<output>
<ID>OUT_1</ID>931 </output>
<output>
<ID>OUT_2</ID>932 </output>
<output>
<ID>OUT_3</ID>933 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>906</ID>
<type>FF_GND</type>
<position>498.5,325</position>
<output>
<ID>OUT_0</ID>934 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>907</ID>
<type>DE_TO</type>
<position>499,278</position>
<input>
<ID>IN_0</ID>991 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 2</lparam></gate>
<gate>
<ID>945</ID>
<type>DE_TO</type>
<position>496,278</position>
<input>
<ID>IN_0</ID>992 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 3</lparam></gate>
<gate>
<ID>946</ID>
<type>DE_TO</type>
<position>533.5,309.5</position>
<input>
<ID>IN_0</ID>932 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>948</ID>
<type>DE_TO</type>
<position>490,277.5</position>
<input>
<ID>IN_0</ID>997 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 4</lparam></gate>
<gate>
<ID>949</ID>
<type>DE_TO</type>
<position>531,309</position>
<input>
<ID>IN_0</ID>931 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>950</ID>
<type>DE_TO</type>
<position>528,309.5</position>
<input>
<ID>IN_0</ID>930 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>951</ID>
<type>DE_TO</type>
<position>524.5,309.5</position>
<input>
<ID>IN_0</ID>929 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>952</ID>
<type>DE_TO</type>
<position>485.5,277.5</position>
<input>
<ID>IN_0</ID>998 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 5</lparam></gate>
<gate>
<ID>953</ID>
<type>DE_TO</type>
<position>522,309.5</position>
<input>
<ID>IN_0</ID>928 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>954</ID>
<type>DE_TO</type>
<position>482.5,277.5</position>
<input>
<ID>IN_0</ID>999 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 6</lparam></gate>
<gate>
<ID>955</ID>
<type>DA_FROM</type>
<position>421,333.5</position>
<input>
<ID>IN_0</ID>949 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>956</ID>
<type>DA_FROM</type>
<position>421,330.5</position>
<input>
<ID>IN_0</ID>950 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>957</ID>
<type>DA_FROM</type>
<position>421,328</position>
<input>
<ID>IN_0</ID>951 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>958</ID>
<type>AI_REGISTER12</type>
<position>458,317.5</position>
<input>
<ID>IN_0</ID>942 </input>
<input>
<ID>IN_1</ID>937 </input>
<input>
<ID>IN_10</ID>946 </input>
<input>
<ID>IN_11</ID>945 </input>
<input>
<ID>IN_2</ID>938 </input>
<input>
<ID>IN_3</ID>939 </input>
<input>
<ID>IN_4</ID>940 </input>
<input>
<ID>IN_5</ID>941 </input>
<input>
<ID>IN_6</ID>936 </input>
<input>
<ID>IN_7</ID>935 </input>
<input>
<ID>IN_8</ID>944 </input>
<input>
<ID>IN_9</ID>943 </input>
<output>
<ID>OUT_0</ID>790 </output>
<output>
<ID>OUT_1</ID>789 </output>
<output>
<ID>OUT_10</ID>769 </output>
<output>
<ID>OUT_11</ID>768 </output>
<output>
<ID>OUT_2</ID>788 </output>
<output>
<ID>OUT_3</ID>791 </output>
<output>
<ID>OUT_4</ID>787 </output>
<output>
<ID>OUT_5</ID>770 </output>
<output>
<ID>OUT_6</ID>767 </output>
<output>
<ID>OUT_7</ID>772 </output>
<output>
<ID>OUT_8</ID>771 </output>
<output>
<ID>OUT_9</ID>766 </output>
<input>
<ID>clear</ID>762 </input>
<input>
<ID>clock</ID>761 </input>
<input>
<ID>count_enable</ID>765 </input>
<input>
<ID>count_up</ID>1003 </input>
<input>
<ID>load</ID>764 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>959</ID>
<type>DA_FROM</type>
<position>421,325.5</position>
<input>
<ID>IN_0</ID>952 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>960</ID>
<type>DE_TO</type>
<position>479,278</position>
<input>
<ID>IN_0</ID>1000 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 7</lparam></gate>
<gate>
<ID>962</ID>
<type>DE_TO</type>
<position>519,309.5</position>
<input>
<ID>IN_0</ID>927 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>963</ID>
<type>DE_TO</type>
<position>516.5,309.5</position>
<input>
<ID>IN_0</ID>926 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>964</ID>
<type>DE_TO</type>
<position>475.5,279</position>
<input>
<ID>IN_0</ID>996 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 8</lparam></gate>
<wire>
<ID>965</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>419.5,283,419.5,288.5</points>
<intersection>283 1</intersection>
<intersection>288.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>419.5,283,425,283</points>
<connection>
<GID>801</GID>
<name>IN_0</name></connection>
<intersection>419.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>414.5,288.5,419.5,288.5</points>
<connection>
<GID>872</GID>
<name>IN_0</name></connection>
<intersection>419.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>772</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>463,319,493.5,319</points>
<connection>
<GID>958</GID>
<name>OUT_7</name></connection>
<connection>
<GID>972</GID>
<name>IN_3</name></connection>
<intersection>480 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>480,296,480,319</points>
<connection>
<GID>986</GID>
<name>IN_3</name></connection>
<intersection>319 1</intersection></vsegment></shape></wire>
<wire>
<ID>966</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>420,272,420,277</points>
<intersection>272 3</intersection>
<intersection>277 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>420,277,429.5,277</points>
<connection>
<GID>799</GID>
<name>IN_2</name></connection>
<intersection>420 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>414.5,272,420,272</points>
<connection>
<GID>680</GID>
<name>IN_0</name></connection>
<intersection>420 0</intersection></hsegment></shape></wire>
<wire>
<ID>967</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>419,275,419,278</points>
<intersection>275 2</intersection>
<intersection>278 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>419,278,429.5,278</points>
<connection>
<GID>799</GID>
<name>IN_3</name></connection>
<intersection>419 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>414.5,275,419,275</points>
<connection>
<GID>898</GID>
<name>IN_0</name></connection>
<intersection>419 0</intersection></hsegment></shape></wire>
<wire>
<ID>968</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>417.5,277.5,417.5,279</points>
<intersection>277.5 1</intersection>
<intersection>279 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>414.5,277.5,417.5,277.5</points>
<connection>
<GID>897</GID>
<name>IN_0</name></connection>
<intersection>417.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>417.5,279,429.5,279</points>
<connection>
<GID>799</GID>
<name>IN_4</name></connection>
<intersection>417.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>969</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>414.5,280,429.5,280</points>
<connection>
<GID>896</GID>
<name>IN_0</name></connection>
<connection>
<GID>799</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>970</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>417.5,281,417.5,283</points>
<intersection>281 2</intersection>
<intersection>283 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>414.5,283,417.5,283</points>
<connection>
<GID>874</GID>
<name>IN_0</name></connection>
<intersection>417.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>417.5,281,429.5,281</points>
<connection>
<GID>799</GID>
<name>IN_6</name></connection>
<intersection>417.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>971</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>419,282,419,285.5</points>
<intersection>282 2</intersection>
<intersection>285.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>414.5,285.5,419,285.5</points>
<connection>
<GID>873</GID>
<name>IN_0</name></connection>
<intersection>419 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>419,282,429.5,282</points>
<connection>
<GID>799</GID>
<name>IN_7</name></connection>
<intersection>419 0</intersection></hsegment></shape></wire>
<wire>
<ID>972</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>427,289.5,431.5,289.5</points>
<connection>
<GID>822</GID>
<name>IN_0</name></connection>
<intersection>427 5</intersection>
<intersection>431.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>431.5,283.5,431.5,289.5</points>
<connection>
<GID>799</GID>
<name>ENABLE_0</name></connection>
<intersection>289.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>427,287.5,427,289.5</points>
<connection>
<GID>801</GID>
<name>ENABLE_0</name></connection>
<intersection>289.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>973</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>493,293,493.5,293</points>
<connection>
<GID>986</GID>
<name>carry_in</name></connection>
<connection>
<GID>988</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>974</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>476.5,293,477,293</points>
<connection>
<GID>984</GID>
<name>carry_in</name></connection>
<connection>
<GID>986</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>975</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510.5,292,510.5,293</points>
<connection>
<GID>990</GID>
<name>OUT_0</name></connection>
<intersection>293 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>509.5,293,510.5,293</points>
<connection>
<GID>988</GID>
<name>carry_in</name></connection>
<intersection>510.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>976</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>503,287,503,288</points>
<connection>
<GID>988</GID>
<name>OUT_0</name></connection>
<connection>
<GID>992</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>977</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502,287,502,288</points>
<connection>
<GID>988</GID>
<name>OUT_1</name></connection>
<connection>
<GID>992</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>978</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>501,287,501,288</points>
<connection>
<GID>988</GID>
<name>OUT_2</name></connection>
<connection>
<GID>992</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>979</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>500,287,500,288</points>
<connection>
<GID>988</GID>
<name>OUT_3</name></connection>
<connection>
<GID>992</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>980</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>483.5,287,483.5,288</points>
<connection>
<GID>986</GID>
<name>OUT_3</name></connection>
<connection>
<GID>994</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>787</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>463,316,493.5,316</points>
<connection>
<GID>958</GID>
<name>OUT_4</name></connection>
<connection>
<GID>972</GID>
<name>IN_0</name></connection>
<intersection>483 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>483,296,483,316</points>
<connection>
<GID>986</GID>
<name>IN_0</name></connection>
<intersection>316 1</intersection></vsegment></shape></wire>
<wire>
<ID>981</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484.5,287,484.5,288</points>
<connection>
<GID>986</GID>
<name>OUT_2</name></connection>
<connection>
<GID>994</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>788</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>463,314,489,314</points>
<connection>
<GID>958</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1</GID>
<name>IN_2</name></connection>
<intersection>486 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>486,299,486,314</points>
<intersection>299 9</intersection>
<intersection>314 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>486,299,497.5,299</points>
<intersection>486 8</intersection>
<intersection>497.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>497.5,296,497.5,299</points>
<connection>
<GID>988</GID>
<name>IN_2</name></connection>
<intersection>299 9</intersection></vsegment></shape></wire>
<wire>
<ID>982</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>486.5,287,486.5,288</points>
<connection>
<GID>986</GID>
<name>OUT_0</name></connection>
<connection>
<GID>994</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>789</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>463,313,489,313</points>
<connection>
<GID>958</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>487.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>487.5,300,487.5,313</points>
<intersection>300 9</intersection>
<intersection>313 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>487.5,300,498.5,300</points>
<intersection>487.5 8</intersection>
<intersection>498.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>498.5,296,498.5,300</points>
<connection>
<GID>988</GID>
<name>IN_1</name></connection>
<intersection>300 9</intersection></vsegment></shape></wire>
<wire>
<ID>983</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>485.5,287,485.5,288</points>
<connection>
<GID>986</GID>
<name>OUT_1</name></connection>
<connection>
<GID>994</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>790</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>463,312,489,312</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<connection>
<GID>958</GID>
<name>OUT_0</name></connection>
<intersection>489 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>489,301,489,312</points>
<intersection>301 9</intersection>
<intersection>312 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>489,301,499.5,301</points>
<intersection>489 8</intersection>
<intersection>499.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>499.5,296,499.5,301</points>
<connection>
<GID>988</GID>
<name>IN_0</name></connection>
<intersection>301 9</intersection></vsegment></shape></wire>
<wire>
<ID>984</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>470,287,470,288</points>
<connection>
<GID>984</GID>
<name>OUT_0</name></connection>
<connection>
<GID>996</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>791</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>463,315,489,315</points>
<connection>
<GID>958</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1</GID>
<name>IN_3</name></connection>
<intersection>485 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>485,297.5,485,315</points>
<intersection>297.5 9</intersection>
<intersection>315 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>485,297.5,496.5,297.5</points>
<intersection>485 8</intersection>
<intersection>496.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>496.5,296,496.5,297.5</points>
<connection>
<GID>988</GID>
<name>IN_3</name></connection>
<intersection>297.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>985</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467,287,467,288</points>
<connection>
<GID>984</GID>
<name>OUT_3</name></connection>
<connection>
<GID>996</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>986</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>469,287,469,288</points>
<connection>
<GID>984</GID>
<name>OUT_1</name></connection>
<connection>
<GID>996</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>987</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>468,287,468,288</points>
<connection>
<GID>984</GID>
<name>OUT_2</name></connection>
<connection>
<GID>996</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>988</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>471.5,285,508,285</points>
<connection>
<GID>996</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>994</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>992</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>659</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>989</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>505,280.5,505,283</points>
<connection>
<GID>901</GID>
<name>IN_0</name></connection>
<intersection>283 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>503,283,505,283</points>
<connection>
<GID>992</GID>
<name>OUT_3</name></connection>
<intersection>505 0</intersection></hsegment></shape></wire>
<wire>
<ID>990</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>502,280,502,283</points>
<connection>
<GID>992</GID>
<name>OUT_2</name></connection>
<connection>
<GID>904</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>991</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>501,281.5,501,283</points>
<connection>
<GID>992</GID>
<name>OUT_1</name></connection>
<intersection>281.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>499,280,499,281.5</points>
<connection>
<GID>907</GID>
<name>IN_0</name></connection>
<intersection>281.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>499,281.5,501,281.5</points>
<intersection>499 1</intersection>
<intersection>501 0</intersection></hsegment></shape></wire>
<wire>
<ID>992</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>500,282,500,283</points>
<connection>
<GID>992</GID>
<name>OUT_0</name></connection>
<intersection>282 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>496,280,496,282</points>
<connection>
<GID>945</GID>
<name>IN_0</name></connection>
<intersection>282 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>496,282,500,282</points>
<intersection>496 1</intersection>
<intersection>500 0</intersection></hsegment></shape></wire>
<wire>
<ID>993</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467,282,467,283</points>
<connection>
<GID>996</GID>
<name>OUT_0</name></connection>
<intersection>282 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>465,280.5,465,282</points>
<connection>
<GID>980</GID>
<name>IN_0</name></connection>
<intersection>282 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>465,282,467,282</points>
<intersection>465 1</intersection>
<intersection>467 0</intersection></hsegment></shape></wire>
<wire>
<ID>994</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>468,280.5,468,283</points>
<connection>
<GID>976</GID>
<name>IN_0</name></connection>
<connection>
<GID>996</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>995</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>469,281.5,469,283</points>
<connection>
<GID>996</GID>
<name>OUT_2</name></connection>
<intersection>281.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>471.5,280.5,471.5,281.5</points>
<connection>
<GID>974</GID>
<name>IN_0</name></connection>
<intersection>281.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>469,281.5,471.5,281.5</points>
<intersection>469 0</intersection>
<intersection>471.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>996</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>470,282,470,283</points>
<connection>
<GID>996</GID>
<name>OUT_3</name></connection>
<intersection>282 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>475.5,281,475.5,282</points>
<connection>
<GID>964</GID>
<name>IN_0</name></connection>
<intersection>282 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>470,282,475.5,282</points>
<intersection>470 0</intersection>
<intersection>475.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>997</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>490,279.5,490,283</points>
<connection>
<GID>948</GID>
<name>IN_0</name></connection>
<intersection>283 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>486.5,283,490,283</points>
<connection>
<GID>994</GID>
<name>OUT_3</name></connection>
<intersection>490 0</intersection></hsegment></shape></wire>
<wire>
<ID>998</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>485.5,279.5,485.5,283</points>
<connection>
<GID>994</GID>
<name>OUT_2</name></connection>
<connection>
<GID>952</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>999</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484.5,281,484.5,283</points>
<connection>
<GID>994</GID>
<name>OUT_1</name></connection>
<intersection>281 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>482.5,279.5,482.5,281</points>
<connection>
<GID>954</GID>
<name>IN_0</name></connection>
<intersection>281 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>482.5,281,484.5,281</points>
<intersection>482.5 1</intersection>
<intersection>484.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1000</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>483.5,281.5,483.5,283</points>
<connection>
<GID>994</GID>
<name>OUT_0</name></connection>
<intersection>281.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>479,280,479,281.5</points>
<connection>
<GID>960</GID>
<name>IN_0</name></connection>
<intersection>281.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>479,281.5,483.5,281.5</points>
<intersection>479 1</intersection>
<intersection>483.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1001</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>506.5,296,506.5,296.5</points>
<connection>
<GID>988</GID>
<name>IN_B_0</name></connection>
<intersection>296.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>470.5,296.5,514,296.5</points>
<connection>
<GID>998</GID>
<name>IN_0</name></connection>
<intersection>470.5 16</intersection>
<intersection>471.5 17</intersection>
<intersection>472.5 18</intersection>
<intersection>473.5 19</intersection>
<intersection>487 20</intersection>
<intersection>488 21</intersection>
<intersection>489 22</intersection>
<intersection>490 23</intersection>
<intersection>503.5 5</intersection>
<intersection>504.5 6</intersection>
<intersection>505.5 7</intersection>
<intersection>506.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>503.5,296,503.5,296.5</points>
<connection>
<GID>988</GID>
<name>IN_B_3</name></connection>
<intersection>296.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>504.5,296,504.5,296.5</points>
<connection>
<GID>988</GID>
<name>IN_B_2</name></connection>
<intersection>296.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>505.5,296,505.5,296.5</points>
<connection>
<GID>988</GID>
<name>IN_B_1</name></connection>
<intersection>296.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>470.5,296,470.5,296.5</points>
<connection>
<GID>984</GID>
<name>IN_B_3</name></connection>
<intersection>296.5 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>471.5,296,471.5,296.5</points>
<connection>
<GID>984</GID>
<name>IN_B_2</name></connection>
<intersection>296.5 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>472.5,296,472.5,296.5</points>
<connection>
<GID>984</GID>
<name>IN_B_1</name></connection>
<intersection>296.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>473.5,296,473.5,296.5</points>
<connection>
<GID>984</GID>
<name>IN_B_0</name></connection>
<intersection>296.5 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>487,296,487,296.5</points>
<connection>
<GID>986</GID>
<name>IN_B_3</name></connection>
<intersection>296.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>488,296,488,296.5</points>
<connection>
<GID>986</GID>
<name>IN_B_2</name></connection>
<intersection>296.5 1</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>489,296,489,296.5</points>
<connection>
<GID>986</GID>
<name>IN_B_1</name></connection>
<intersection>296.5 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>490,296,490,296.5</points>
<connection>
<GID>986</GID>
<name>IN_B_0</name></connection>
<intersection>296.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1002</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>469.5,327.5,469.5,327.5</points>
<connection>
<GID>999</GID>
<name>IN_0</name></connection>
<connection>
<GID>1001</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1003</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459,325,459,327.5</points>
<connection>
<GID>958</GID>
<name>count_up</name></connection>
<intersection>327.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>459,327.5,465.5,327.5</points>
<connection>
<GID>1001</GID>
<name>OUT_0</name></connection>
<intersection>459 0</intersection></hsegment></shape></wire>
<wire>
<ID>870</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491,316.5,491,331.5</points>
<connection>
<GID>1</GID>
<name>ENABLE_0</name></connection>
<intersection>324.5 13</intersection>
<intersection>331.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>491,331.5,501.5,331.5</points>
<connection>
<GID>905</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>899</GID>
<name>IN_0</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>491,324.5,495.5,324.5</points>
<connection>
<GID>972</GID>
<name>ENABLE_0</name></connection>
<intersection>491 0</intersection></hsegment></shape></wire>
<wire>
<ID>918</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>493,312,494,312</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>494 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>494,311,494,312</points>
<connection>
<GID>965</GID>
<name>IN_0</name></connection>
<intersection>312 1</intersection></vsegment></shape></wire>
<wire>
<ID>919</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497.5,311,497.5,313</points>
<connection>
<GID>966</GID>
<name>IN_0</name></connection>
<intersection>313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>493,313,497.5,313</points>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection>
<intersection>497.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>920</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>500.5,311,500.5,314</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>314 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>493,314,500.5,314</points>
<connection>
<GID>1</GID>
<name>OUT_2</name></connection>
<intersection>500.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>921</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>503.5,311,503.5,315</points>
<connection>
<GID>676</GID>
<name>IN_0</name></connection>
<intersection>315 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>493,315,503.5,315</points>
<connection>
<GID>1</GID>
<name>OUT_3</name></connection>
<intersection>503.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>922</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>506.5,311,506.5,316</points>
<connection>
<GID>682</GID>
<name>IN_0</name></connection>
<intersection>316 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>497.5,316,506.5,316</points>
<connection>
<GID>972</GID>
<name>OUT_0</name></connection>
<intersection>506.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>923</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>509,311,509,317</points>
<connection>
<GID>885</GID>
<name>IN_0</name></connection>
<intersection>317 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>497.5,317,509,317</points>
<connection>
<GID>972</GID>
<name>OUT_1</name></connection>
<intersection>509 0</intersection></hsegment></shape></wire>
<wire>
<ID>924</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511.5,311.5,511.5,318</points>
<connection>
<GID>902</GID>
<name>IN_0</name></connection>
<intersection>318 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>497.5,318,511.5,318</points>
<connection>
<GID>972</GID>
<name>OUT_2</name></connection>
<intersection>511.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>925</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513.5,311.5,513.5,319</points>
<connection>
<GID>903</GID>
<name>IN_0</name></connection>
<intersection>319 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>497.5,319,513.5,319</points>
<connection>
<GID>972</GID>
<name>OUT_3</name></connection>
<intersection>513.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>926</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516.5,311.5,516.5,320</points>
<connection>
<GID>963</GID>
<name>IN_0</name></connection>
<intersection>320 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>497.5,320,516.5,320</points>
<connection>
<GID>972</GID>
<name>OUT_4</name></connection>
<intersection>516.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>927</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>519,311.5,519,321</points>
<connection>
<GID>962</GID>
<name>IN_0</name></connection>
<intersection>321 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>497.5,321,519,321</points>
<connection>
<GID>972</GID>
<name>OUT_5</name></connection>
<intersection>519 0</intersection></hsegment></shape></wire>
<wire>
<ID>928</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>522,311.5,522,322</points>
<connection>
<GID>953</GID>
<name>IN_0</name></connection>
<intersection>322 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>497.5,322,522,322</points>
<connection>
<GID>972</GID>
<name>OUT_6</name></connection>
<intersection>522 0</intersection></hsegment></shape></wire>
<wire>
<ID>929</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>524.5,311.5,524.5,323</points>
<connection>
<GID>951</GID>
<name>IN_0</name></connection>
<intersection>323 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>497.5,323,524.5,323</points>
<connection>
<GID>972</GID>
<name>OUT_7</name></connection>
<intersection>524.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>930</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>528,311.5,528,327</points>
<connection>
<GID>950</GID>
<name>IN_0</name></connection>
<intersection>327 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>503.5,327,528,327</points>
<connection>
<GID>905</GID>
<name>OUT_0</name></connection>
<intersection>528 0</intersection></hsegment></shape></wire>
<wire>
<ID>931</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>531,311,531,328</points>
<connection>
<GID>949</GID>
<name>IN_0</name></connection>
<intersection>328 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>503.5,328,531,328</points>
<connection>
<GID>905</GID>
<name>OUT_1</name></connection>
<intersection>531 0</intersection></hsegment></shape></wire>
<wire>
<ID>932</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>533.5,311.5,533.5,329</points>
<connection>
<GID>946</GID>
<name>IN_0</name></connection>
<intersection>329 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>503.5,329,533.5,329</points>
<connection>
<GID>905</GID>
<name>OUT_2</name></connection>
<intersection>533.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>933</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>536.5,311,536.5,330</points>
<connection>
<GID>663</GID>
<name>IN_0</name></connection>
<intersection>330 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>503.5,330,536.5,330</points>
<connection>
<GID>905</GID>
<name>OUT_3</name></connection>
<intersection>536.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>934</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>498.5,326,498.5,327</points>
<connection>
<GID>906</GID>
<name>OUT_0</name></connection>
<intersection>327 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>498.5,327,499.5,327</points>
<connection>
<GID>905</GID>
<name>IN_0</name></connection>
<intersection>498.5 0</intersection>
<intersection>499.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>499.5,327,499.5,330</points>
<connection>
<GID>905</GID>
<name>IN_3</name></connection>
<connection>
<GID>905</GID>
<name>IN_2</name></connection>
<connection>
<GID>905</GID>
<name>IN_1</name></connection>
<intersection>327 1</intersection></vsegment></shape></wire>
<wire>
<ID>935</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440.5,319,453,319</points>
<connection>
<GID>958</GID>
<name>IN_7</name></connection>
<connection>
<GID>661</GID>
<name>OUT_7</name></connection>
<intersection>446 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>446,282,446,319</points>
<intersection>282 7</intersection>
<intersection>319 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>433.5,282,446,282</points>
<connection>
<GID>799</GID>
<name>OUT_7</name></connection>
<intersection>446 6</intersection></hsegment></shape></wire>
<wire>
<ID>936</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440.5,318,453,318</points>
<connection>
<GID>958</GID>
<name>IN_6</name></connection>
<connection>
<GID>661</GID>
<name>OUT_6</name></connection>
<intersection>447 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>447,281,447,318</points>
<intersection>281 7</intersection>
<intersection>318 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>433.5,281,447,281</points>
<connection>
<GID>799</GID>
<name>OUT_6</name></connection>
<intersection>447 6</intersection></hsegment></shape></wire>
<wire>
<ID>937</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440.5,313,453,313</points>
<connection>
<GID>958</GID>
<name>IN_1</name></connection>
<connection>
<GID>661</GID>
<name>OUT_1</name></connection>
<intersection>452 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>452,276,452,313</points>
<intersection>276 16</intersection>
<intersection>313 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>433.5,276,452,276</points>
<connection>
<GID>799</GID>
<name>OUT_1</name></connection>
<intersection>452 15</intersection></hsegment></shape></wire>
<wire>
<ID>938</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440.5,314,453,314</points>
<connection>
<GID>958</GID>
<name>IN_2</name></connection>
<connection>
<GID>661</GID>
<name>OUT_2</name></connection>
<intersection>451 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>451,277,451,314</points>
<intersection>277 16</intersection>
<intersection>314 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>433.5,277,451,277</points>
<connection>
<GID>799</GID>
<name>OUT_2</name></connection>
<intersection>451 15</intersection></hsegment></shape></wire>
<wire>
<ID>939</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440.5,315,453,315</points>
<connection>
<GID>958</GID>
<name>IN_3</name></connection>
<connection>
<GID>661</GID>
<name>OUT_3</name></connection>
<intersection>450 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>450,278,450,315</points>
<intersection>278 16</intersection>
<intersection>315 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>433.5,278,450,278</points>
<connection>
<GID>799</GID>
<name>OUT_3</name></connection>
<intersection>450 15</intersection></hsegment></shape></wire>
<wire>
<ID>940</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440.5,316,453,316</points>
<connection>
<GID>958</GID>
<name>IN_4</name></connection>
<connection>
<GID>661</GID>
<name>OUT_4</name></connection>
<intersection>449 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>449,279,449,316</points>
<intersection>279 10</intersection>
<intersection>316 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>433.5,279,449,279</points>
<connection>
<GID>799</GID>
<name>OUT_4</name></connection>
<intersection>449 9</intersection></hsegment></shape></wire>
<wire>
<ID>941</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440.5,317,453,317</points>
<connection>
<GID>958</GID>
<name>IN_5</name></connection>
<connection>
<GID>661</GID>
<name>OUT_5</name></connection>
<intersection>448 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>448,280,448,317</points>
<intersection>280 10</intersection>
<intersection>317 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>433.5,280,448,280</points>
<connection>
<GID>799</GID>
<name>OUT_5</name></connection>
<intersection>448 9</intersection></hsegment></shape></wire>
<wire>
<ID>942</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>440.5,312,453,312</points>
<connection>
<GID>958</GID>
<name>IN_0</name></connection>
<connection>
<GID>661</GID>
<name>OUT_0</name></connection>
<intersection>453 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>453,275,453,312</points>
<intersection>275 16</intersection>
<intersection>312 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>433.5,275,453,275</points>
<connection>
<GID>799</GID>
<name>OUT_0</name></connection>
<intersection>453 15</intersection></hsegment></shape></wire>
<wire>
<ID>943</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>436.5,321,453,321</points>
<connection>
<GID>958</GID>
<name>IN_9</name></connection>
<connection>
<GID>667</GID>
<name>OUT_1</name></connection>
<intersection>444 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>444,284,444,321</points>
<intersection>284 7</intersection>
<intersection>321 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>429,284,444,284</points>
<connection>
<GID>801</GID>
<name>OUT_1</name></connection>
<intersection>444 6</intersection></hsegment></shape></wire>
<wire>
<ID>944</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>436.5,320,453,320</points>
<connection>
<GID>958</GID>
<name>IN_8</name></connection>
<connection>
<GID>667</GID>
<name>OUT_0</name></connection>
<intersection>445 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>445,283,445,320</points>
<intersection>283 7</intersection>
<intersection>320 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>429,283,445,283</points>
<connection>
<GID>801</GID>
<name>OUT_0</name></connection>
<intersection>445 6</intersection></hsegment></shape></wire>
<wire>
<ID>945</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>436.5,323,453,323</points>
<connection>
<GID>958</GID>
<name>IN_11</name></connection>
<connection>
<GID>667</GID>
<name>OUT_3</name></connection>
<intersection>442 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>442,286,442,323</points>
<intersection>286 7</intersection>
<intersection>323 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>429,286,442,286</points>
<connection>
<GID>801</GID>
<name>OUT_3</name></connection>
<intersection>442 6</intersection></hsegment></shape></wire>
<wire>
<ID>946</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>436.5,322,453,322</points>
<connection>
<GID>958</GID>
<name>IN_10</name></connection>
<connection>
<GID>667</GID>
<name>OUT_2</name></connection>
<intersection>443 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>443,285,443,322</points>
<intersection>285 7</intersection>
<intersection>322 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>429,285,443,285</points>
<connection>
<GID>801</GID>
<name>OUT_2</name></connection>
<intersection>443 6</intersection></hsegment></shape></wire>
<wire>
<ID>947</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431,303,431,312</points>
<intersection>303 2</intersection>
<intersection>312 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>422.5,303,431,303</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>431 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>431,312,436.5,312</points>
<connection>
<GID>661</GID>
<name>IN_0</name></connection>
<intersection>431 0</intersection></hsegment></shape></wire>
<wire>
<ID>948</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430,306,430,313</points>
<intersection>306 2</intersection>
<intersection>313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>430,313,436.5,313</points>
<connection>
<GID>661</GID>
<name>IN_1</name></connection>
<intersection>430 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>422.5,306,430,306</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>430 0</intersection></hsegment></shape></wire>
<wire>
<ID>949</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432,323,432,333.5</points>
<intersection>323 2</intersection>
<intersection>333.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423,333.5,432,333.5</points>
<connection>
<GID>955</GID>
<name>IN_0</name></connection>
<intersection>432 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>432,323,432.5,323</points>
<connection>
<GID>667</GID>
<name>IN_3</name></connection>
<intersection>432 0</intersection></hsegment></shape></wire>
<wire>
<ID>950</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430.5,322,430.5,330.5</points>
<intersection>322 2</intersection>
<intersection>330.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423,330.5,430.5,330.5</points>
<connection>
<GID>956</GID>
<name>IN_0</name></connection>
<intersection>430.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>430.5,322,432.5,322</points>
<connection>
<GID>667</GID>
<name>IN_2</name></connection>
<intersection>430.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>951</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429.5,321,429.5,328</points>
<intersection>321 3</intersection>
<intersection>328 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>423,328,429.5,328</points>
<connection>
<GID>957</GID>
<name>IN_0</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>429.5,321,432.5,321</points>
<connection>
<GID>667</GID>
<name>IN_1</name></connection>
<intersection>429.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>952</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428,320,428,325.5</points>
<intersection>320 1</intersection>
<intersection>325.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428,320,432.5,320</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>428 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>423,325.5,428,325.5</points>
<connection>
<GID>959</GID>
<name>IN_0</name></connection>
<intersection>428 0</intersection></hsegment></shape></wire>
<wire>
<ID>953</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428.5,309,428.5,314</points>
<intersection>309 3</intersection>
<intersection>314 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,314,436.5,314</points>
<connection>
<GID>661</GID>
<name>IN_2</name></connection>
<intersection>428.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>423,309,428.5,309</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>428.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>954</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,312,427.5,315</points>
<intersection>312 2</intersection>
<intersection>315 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427.5,315,436.5,315</points>
<connection>
<GID>661</GID>
<name>IN_3</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>423,312,427.5,312</points>
<connection>
<GID>979</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>761</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457,308,457,310</points>
<connection>
<GID>958</GID>
<name>clock</name></connection>
<connection>
<GID>967</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>955</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426,314.5,426,316</points>
<intersection>314.5 1</intersection>
<intersection>316 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423,314.5,426,314.5</points>
<connection>
<GID>978</GID>
<name>IN_0</name></connection>
<intersection>426 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>426,316,436.5,316</points>
<connection>
<GID>661</GID>
<name>IN_4</name></connection>
<intersection>426 0</intersection></hsegment></shape></wire>
<wire>
<ID>762</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>459,308.5,459,310</points>
<connection>
<GID>958</GID>
<name>clear</name></connection>
<connection>
<GID>968</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>956</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>423,317,436.5,317</points>
<connection>
<GID>661</GID>
<name>IN_5</name></connection>
<connection>
<GID>977</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>957</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426,318,426,320</points>
<intersection>318 2</intersection>
<intersection>320 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423,320,426,320</points>
<connection>
<GID>975</GID>
<name>IN_0</name></connection>
<intersection>426 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>426,318,436.5,318</points>
<connection>
<GID>661</GID>
<name>IN_6</name></connection>
<intersection>426 0</intersection></hsegment></shape></wire>
<wire>
<ID>764</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>457,325,457,333.5</points>
<connection>
<GID>958</GID>
<name>load</name></connection>
<intersection>333.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>453,333.5,457,333.5</points>
<connection>
<GID>970</GID>
<name>IN_0</name></connection>
<intersection>457 0</intersection></hsegment></shape></wire>
<wire>
<ID>958</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,319,427.5,322.5</points>
<intersection>319 2</intersection>
<intersection>322.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423,322.5,427.5,322.5</points>
<connection>
<GID>973</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>427.5,319,436.5,319</points>
<connection>
<GID>661</GID>
<name>IN_7</name></connection>
<intersection>427.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>765</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458,325,458,337</points>
<connection>
<GID>958</GID>
<name>count_enable</name></connection>
<intersection>337 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>452,337,458,337</points>
<connection>
<GID>971</GID>
<name>IN_0</name></connection>
<intersection>458 0</intersection></hsegment></shape></wire>
<wire>
<ID>959</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,324.5,434.5,328</points>
<connection>
<GID>667</GID>
<name>ENABLE_0</name></connection>
<intersection>324.5 2</intersection>
<intersection>328 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434.5,328,437.5,328</points>
<connection>
<GID>678</GID>
<name>IN_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>434.5,324.5,438.5,324.5</points>
<intersection>434.5 0</intersection>
<intersection>438.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>438.5,320.5,438.5,324.5</points>
<connection>
<GID>661</GID>
<name>ENABLE_0</name></connection>
<intersection>324.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>766</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>463,321,493.5,321</points>
<connection>
<GID>958</GID>
<name>OUT_9</name></connection>
<connection>
<GID>972</GID>
<name>IN_5</name></connection>
<intersection>465.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>465.5,296,465.5,321</points>
<connection>
<GID>984</GID>
<name>IN_1</name></connection>
<intersection>321 1</intersection></vsegment></shape></wire>
<wire>
<ID>960</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>422.5,266,422.5,275</points>
<intersection>266 2</intersection>
<intersection>275 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>414,266,422.5,266</points>
<connection>
<GID>797</GID>
<name>IN_0</name></connection>
<intersection>422.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>422.5,275,429.5,275</points>
<connection>
<GID>799</GID>
<name>IN_0</name></connection>
<intersection>422.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>767</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>463,318,493.5,318</points>
<connection>
<GID>958</GID>
<name>OUT_6</name></connection>
<connection>
<GID>972</GID>
<name>IN_2</name></connection>
<intersection>481 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>481,296,481,318</points>
<connection>
<GID>986</GID>
<name>IN_2</name></connection>
<intersection>318 1</intersection></vsegment></shape></wire>
<wire>
<ID>961</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421.5,269,421.5,276</points>
<intersection>269 2</intersection>
<intersection>276 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>421.5,276,429.5,276</points>
<connection>
<GID>799</GID>
<name>IN_1</name></connection>
<intersection>421.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>414,269,421.5,269</points>
<connection>
<GID>684</GID>
<name>IN_0</name></connection>
<intersection>421.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>768</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>463,323,493.5,323</points>
<connection>
<GID>958</GID>
<name>OUT_11</name></connection>
<connection>
<GID>972</GID>
<name>IN_7</name></connection>
<intersection>463.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>463.5,296,463.5,323</points>
<connection>
<GID>984</GID>
<name>IN_3</name></connection>
<intersection>323 1</intersection></vsegment></shape></wire>
<wire>
<ID>962</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>423.5,286,423.5,296.5</points>
<intersection>286 2</intersection>
<intersection>296.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>414.5,296.5,423.5,296.5</points>
<connection>
<GID>828</GID>
<name>IN_0</name></connection>
<intersection>423.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>423.5,286,425,286</points>
<connection>
<GID>801</GID>
<name>IN_3</name></connection>
<intersection>423.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>769</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>463,322,493.5,322</points>
<connection>
<GID>958</GID>
<name>OUT_10</name></connection>
<connection>
<GID>972</GID>
<name>IN_6</name></connection>
<intersection>464.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>464.5,296,464.5,322</points>
<connection>
<GID>984</GID>
<name>IN_2</name></connection>
<intersection>322 1</intersection></vsegment></shape></wire>
<wire>
<ID>963</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>422,285,422,293.5</points>
<intersection>285 2</intersection>
<intersection>293.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>414.5,293.5,422,293.5</points>
<connection>
<GID>870</GID>
<name>IN_0</name></connection>
<intersection>422 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>422,285,425,285</points>
<connection>
<GID>801</GID>
<name>IN_2</name></connection>
<intersection>422 0</intersection></hsegment></shape></wire>
<wire>
<ID>770</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>463,317,493.5,317</points>
<connection>
<GID>972</GID>
<name>IN_1</name></connection>
<connection>
<GID>958</GID>
<name>OUT_5</name></connection>
<intersection>482 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>482,296,482,317</points>
<connection>
<GID>986</GID>
<name>IN_1</name></connection>
<intersection>317 1</intersection></vsegment></shape></wire>
<wire>
<ID>964</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421,284,421,291</points>
<intersection>284 3</intersection>
<intersection>291 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>414.5,291,421,291</points>
<connection>
<GID>871</GID>
<name>IN_0</name></connection>
<intersection>421 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>421,284,425,284</points>
<connection>
<GID>801</GID>
<name>IN_1</name></connection>
<intersection>421 0</intersection></hsegment></shape></wire>
<wire>
<ID>771</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>463,320,493.5,320</points>
<connection>
<GID>958</GID>
<name>OUT_8</name></connection>
<connection>
<GID>972</GID>
<name>IN_4</name></connection>
<intersection>466.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>466.5,296,466.5,320</points>
<connection>
<GID>984</GID>
<name>IN_0</name></connection>
<intersection>320 1</intersection></vsegment></shape></wire></page 7>
<page 8>
<PageViewport>-0.001945,1359.91,1126,713.91</PageViewport></page 8>
<page 9>
<PageViewport>-405.916,1626.85,720.084,980.853</PageViewport>
<gate>
<ID>1075</ID>
<type>AA_LABEL</type>
<position>110,1316</position>
<gparam>LABEL_TEXT plagiarism</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate></page 9></circuit>